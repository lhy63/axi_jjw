// Generator : SpinalHDL v1.5.0    git head : 83a031922866b078c411ec5529e00f1b6e79f8e7
// Component : TopAxiMasterWandRWithSlave



module TopAxiMasterWandRWithSlave (
  output              io_rdataOut_valid,
  input               io_rdataOut_ready,
  output     [7:0]    io_rdataOut_payload,
  input               io_rapStart,
  input      [31:0]   io_RAddrOffset,
  input      [31:0]   io_Rlen,
  output              io_rapDone,
  input               io_wapStart,
  input               io_wdata_in_valid,
  output              io_wdata_in_ready,
  input      [7:0]    io_wdata_in_payload,
  input      [31:0]   io_WAddrOffset,
  input      [31:0]   io_Wlen,
  output              io_wapDone,
  input               clk,
  input               reset
);
  wire                axiSlave_apstart;
  wire                axiSlave_axiSignal_ar_ready;
  wire                axiSlave_axiSignal_aw_ready;
  wire                axiSlave_axiSignal_w_ready;
  wire                axiSlave_axiSignal_r_valid;
  wire       [7:0]    axiSlave_axiSignal_r_payload_data;
  wire       [3:0]    axiSlave_axiSignal_r_payload_id;
  wire       [1:0]    axiSlave_axiSignal_r_payload_resp;
  wire                axiSlave_axiSignal_r_payload_last;
  wire                axiSlave_axiSignal_b_valid;
  wire       [3:0]    axiSlave_axiSignal_b_payload_id;
  wire       [1:0]    axiSlave_axiSignal_b_payload_resp;
  wire                axiMasterRead_io_dataOut_valid;
  wire       [7:0]    axiMasterRead_io_dataOut_payload;
  wire                axiMasterRead_io_apDone;
  wire                axiMasterRead_io_axiAR_valid;
  wire       [31:0]   axiMasterRead_io_axiAR_payload_addr;
  wire       [3:0]    axiMasterRead_io_axiAR_payload_id;
  wire       [3:0]    axiMasterRead_io_axiAR_payload_region;
  wire       [7:0]    axiMasterRead_io_axiAR_payload_len;
  wire       [2:0]    axiMasterRead_io_axiAR_payload_size;
  wire       [1:0]    axiMasterRead_io_axiAR_payload_burst;
  wire       [0:0]    axiMasterRead_io_axiAR_payload_lock;
  wire       [3:0]    axiMasterRead_io_axiAR_payload_cache;
  wire       [3:0]    axiMasterRead_io_axiAR_payload_qos;
  wire       [0:0]    axiMasterRead_io_axiAR_payload_user;
  wire       [2:0]    axiMasterRead_io_axiAR_payload_prot;
  wire                axiMasterRead_io_axiR_ready;
  wire                axiMasterWrite_io_data_in_ready;
  wire                axiMasterWrite_io_axiAW_valid;
  wire       [31:0]   axiMasterWrite_io_axiAW_payload_addr;
  wire       [3:0]    axiMasterWrite_io_axiAW_payload_id;
  wire       [3:0]    axiMasterWrite_io_axiAW_payload_region;
  wire       [7:0]    axiMasterWrite_io_axiAW_payload_len;
  wire       [2:0]    axiMasterWrite_io_axiAW_payload_size;
  wire       [1:0]    axiMasterWrite_io_axiAW_payload_burst;
  wire       [0:0]    axiMasterWrite_io_axiAW_payload_lock;
  wire       [3:0]    axiMasterWrite_io_axiAW_payload_cache;
  wire       [3:0]    axiMasterWrite_io_axiAW_payload_qos;
  wire       [0:0]    axiMasterWrite_io_axiAW_payload_user;
  wire       [2:0]    axiMasterWrite_io_axiAW_payload_prot;
  wire                axiMasterWrite_io_axiW_valid;
  wire       [7:0]    axiMasterWrite_io_axiW_payload_data;
  wire       [0:0]    axiMasterWrite_io_axiW_payload_strb;
  wire                axiMasterWrite_io_axiW_payload_last;
  wire                axiMasterWrite_io_axiB_ready;
  wire                axiMasterWrite_io_apDone;

  Axi4_transmission axiSlave (
    .axiSignal_aw_valid             (axiMasterWrite_io_axiAW_valid           ), //i
    .axiSignal_aw_ready             (axiSlave_axiSignal_aw_ready             ), //o
    .axiSignal_aw_payload_addr      (axiMasterWrite_io_axiAW_payload_addr    ), //i
    .axiSignal_aw_payload_id        (axiMasterWrite_io_axiAW_payload_id      ), //i
    .axiSignal_aw_payload_region    (axiMasterWrite_io_axiAW_payload_region  ), //i
    .axiSignal_aw_payload_len       (axiMasterWrite_io_axiAW_payload_len     ), //i
    .axiSignal_aw_payload_size      (axiMasterWrite_io_axiAW_payload_size    ), //i
    .axiSignal_aw_payload_burst     (axiMasterWrite_io_axiAW_payload_burst   ), //i
    .axiSignal_aw_payload_lock      (axiMasterWrite_io_axiAW_payload_lock    ), //i
    .axiSignal_aw_payload_cache     (axiMasterWrite_io_axiAW_payload_cache   ), //i
    .axiSignal_aw_payload_qos       (axiMasterWrite_io_axiAW_payload_qos     ), //i
    .axiSignal_aw_payload_user      (axiMasterWrite_io_axiAW_payload_user    ), //i
    .axiSignal_aw_payload_prot      (axiMasterWrite_io_axiAW_payload_prot    ), //i
    .axiSignal_w_valid              (axiMasterWrite_io_axiW_valid            ), //i
    .axiSignal_w_ready              (axiSlave_axiSignal_w_ready              ), //o
    .axiSignal_w_payload_data       (axiMasterWrite_io_axiW_payload_data     ), //i
    .axiSignal_w_payload_strb       (axiMasterWrite_io_axiW_payload_strb     ), //i
    .axiSignal_w_payload_last       (axiMasterWrite_io_axiW_payload_last     ), //i
    .axiSignal_b_valid              (axiSlave_axiSignal_b_valid              ), //o
    .axiSignal_b_ready              (axiMasterWrite_io_axiB_ready            ), //i
    .axiSignal_b_payload_id         (axiSlave_axiSignal_b_payload_id         ), //o
    .axiSignal_b_payload_resp       (axiSlave_axiSignal_b_payload_resp       ), //o
    .axiSignal_ar_valid             (axiMasterRead_io_axiAR_valid            ), //i
    .axiSignal_ar_ready             (axiSlave_axiSignal_ar_ready             ), //o
    .axiSignal_ar_payload_addr      (axiMasterRead_io_axiAR_payload_addr     ), //i
    .axiSignal_ar_payload_id        (axiMasterRead_io_axiAR_payload_id       ), //i
    .axiSignal_ar_payload_region    (axiMasterRead_io_axiAR_payload_region   ), //i
    .axiSignal_ar_payload_len       (axiMasterRead_io_axiAR_payload_len      ), //i
    .axiSignal_ar_payload_size      (axiMasterRead_io_axiAR_payload_size     ), //i
    .axiSignal_ar_payload_burst     (axiMasterRead_io_axiAR_payload_burst    ), //i
    .axiSignal_ar_payload_lock      (axiMasterRead_io_axiAR_payload_lock     ), //i
    .axiSignal_ar_payload_cache     (axiMasterRead_io_axiAR_payload_cache    ), //i
    .axiSignal_ar_payload_qos       (axiMasterRead_io_axiAR_payload_qos      ), //i
    .axiSignal_ar_payload_user      (axiMasterRead_io_axiAR_payload_user     ), //i
    .axiSignal_ar_payload_prot      (axiMasterRead_io_axiAR_payload_prot     ), //i
    .axiSignal_r_valid              (axiSlave_axiSignal_r_valid              ), //o
    .axiSignal_r_ready              (axiMasterRead_io_axiR_ready             ), //i
    .axiSignal_r_payload_data       (axiSlave_axiSignal_r_payload_data       ), //o
    .axiSignal_r_payload_id         (axiSlave_axiSignal_r_payload_id         ), //o
    .axiSignal_r_payload_resp       (axiSlave_axiSignal_r_payload_resp       ), //o
    .axiSignal_r_payload_last       (axiSlave_axiSignal_r_payload_last       ), //o
    .apstart                        (axiSlave_apstart                        ), //i
    .axireset                       (1'b0                                    ), //i
    .clk                            (clk                                     ), //i
    .reset                          (reset                                   )  //i
  );
  AXI4MasterRead axiMasterRead (
    .io_dataOut_valid           (axiMasterRead_io_dataOut_valid         ), //o
    .io_dataOut_ready           (io_rdataOut_ready                      ), //i
    .io_dataOut_payload         (axiMasterRead_io_dataOut_payload       ), //o
    .io_apStart                 (io_rapStart                            ), //i
    .io_RAddrOffset             (io_RAddrOffset                         ), //i
    .io_Rlen                    (io_Rlen                                ), //i
    .io_apDone                  (axiMasterRead_io_apDone                ), //o
    .io_axiAR_valid             (axiMasterRead_io_axiAR_valid           ), //o
    .io_axiAR_ready             (axiSlave_axiSignal_ar_ready            ), //i
    .io_axiAR_payload_addr      (axiMasterRead_io_axiAR_payload_addr    ), //o
    .io_axiAR_payload_id        (axiMasterRead_io_axiAR_payload_id      ), //o
    .io_axiAR_payload_region    (axiMasterRead_io_axiAR_payload_region  ), //o
    .io_axiAR_payload_len       (axiMasterRead_io_axiAR_payload_len     ), //o
    .io_axiAR_payload_size      (axiMasterRead_io_axiAR_payload_size    ), //o
    .io_axiAR_payload_burst     (axiMasterRead_io_axiAR_payload_burst   ), //o
    .io_axiAR_payload_lock      (axiMasterRead_io_axiAR_payload_lock    ), //o
    .io_axiAR_payload_cache     (axiMasterRead_io_axiAR_payload_cache   ), //o
    .io_axiAR_payload_qos       (axiMasterRead_io_axiAR_payload_qos     ), //o
    .io_axiAR_payload_user      (axiMasterRead_io_axiAR_payload_user    ), //o
    .io_axiAR_payload_prot      (axiMasterRead_io_axiAR_payload_prot    ), //o
    .io_axiR_valid              (axiSlave_axiSignal_r_valid             ), //i
    .io_axiR_ready              (axiMasterRead_io_axiR_ready            ), //o
    .io_axiR_payload_data       (axiSlave_axiSignal_r_payload_data      ), //i
    .io_axiR_payload_id         (axiSlave_axiSignal_r_payload_id        ), //i
    .io_axiR_payload_resp       (axiSlave_axiSignal_r_payload_resp      ), //i
    .io_axiR_payload_last       (axiSlave_axiSignal_r_payload_last      ), //i
    .clk                        (clk                                    ), //i
    .reset                      (reset                                  )  //i
  );
  AXI4MasterWriteWithBuffer axiMasterWrite (
    .io_apStart                 (io_wapStart                             ), //i
    .io_data_in_valid           (io_wdata_in_valid                       ), //i
    .io_data_in_ready           (axiMasterWrite_io_data_in_ready         ), //o
    .io_data_in_payload         (io_wdata_in_payload                     ), //i
    .io_WAddrOffset             (io_WAddrOffset                          ), //i
    .io_Wlen                    (io_Wlen                                 ), //i
    .io_axiAW_valid             (axiMasterWrite_io_axiAW_valid           ), //o
    .io_axiAW_ready             (axiSlave_axiSignal_aw_ready             ), //i
    .io_axiAW_payload_addr      (axiMasterWrite_io_axiAW_payload_addr    ), //o
    .io_axiAW_payload_id        (axiMasterWrite_io_axiAW_payload_id      ), //o
    .io_axiAW_payload_region    (axiMasterWrite_io_axiAW_payload_region  ), //o
    .io_axiAW_payload_len       (axiMasterWrite_io_axiAW_payload_len     ), //o
    .io_axiAW_payload_size      (axiMasterWrite_io_axiAW_payload_size    ), //o
    .io_axiAW_payload_burst     (axiMasterWrite_io_axiAW_payload_burst   ), //o
    .io_axiAW_payload_lock      (axiMasterWrite_io_axiAW_payload_lock    ), //o
    .io_axiAW_payload_cache     (axiMasterWrite_io_axiAW_payload_cache   ), //o
    .io_axiAW_payload_qos       (axiMasterWrite_io_axiAW_payload_qos     ), //o
    .io_axiAW_payload_user      (axiMasterWrite_io_axiAW_payload_user    ), //o
    .io_axiAW_payload_prot      (axiMasterWrite_io_axiAW_payload_prot    ), //o
    .io_axiW_valid              (axiMasterWrite_io_axiW_valid            ), //o
    .io_axiW_ready              (axiSlave_axiSignal_w_ready              ), //i
    .io_axiW_payload_data       (axiMasterWrite_io_axiW_payload_data     ), //o
    .io_axiW_payload_strb       (axiMasterWrite_io_axiW_payload_strb     ), //o
    .io_axiW_payload_last       (axiMasterWrite_io_axiW_payload_last     ), //o
    .io_axiB_valid              (axiSlave_axiSignal_b_valid              ), //i
    .io_axiB_ready              (axiMasterWrite_io_axiB_ready            ), //o
    .io_axiB_payload_id         (axiSlave_axiSignal_b_payload_id         ), //i
    .io_axiB_payload_resp       (axiSlave_axiSignal_b_payload_resp       ), //i
    .io_apDone                  (axiMasterWrite_io_apDone                ), //o
    .clk                        (clk                                     ), //i
    .reset                      (reset                                   )  //i
  );
  assign io_rdataOut_valid = axiMasterRead_io_dataOut_valid;
  assign io_rdataOut_payload = axiMasterRead_io_dataOut_payload;
  assign io_rapDone = axiMasterRead_io_apDone;
  assign axiSlave_apstart = (io_wapStart || io_rapStart);
  assign io_wapDone = axiMasterWrite_io_apDone;
  assign io_wdata_in_ready = axiMasterWrite_io_data_in_ready;

endmodule

module AXI4MasterWriteWithBuffer (
  input               io_apStart,
  input               io_data_in_valid,
  output              io_data_in_ready,
  input      [7:0]    io_data_in_payload,
  input      [31:0]   io_WAddrOffset,
  input      [31:0]   io_Wlen,
  output reg          io_axiAW_valid,
  input               io_axiAW_ready,
  output reg [31:0]   io_axiAW_payload_addr,
  output reg [3:0]    io_axiAW_payload_id,
  output reg [3:0]    io_axiAW_payload_region,
  output reg [7:0]    io_axiAW_payload_len,
  output reg [2:0]    io_axiAW_payload_size,
  output reg [1:0]    io_axiAW_payload_burst,
  output reg [0:0]    io_axiAW_payload_lock,
  output reg [3:0]    io_axiAW_payload_cache,
  output reg [3:0]    io_axiAW_payload_qos,
  output reg [0:0]    io_axiAW_payload_user,
  output reg [2:0]    io_axiAW_payload_prot,
  output              io_axiW_valid,
  input               io_axiW_ready,
  output     [7:0]    io_axiW_payload_data,
  output     [0:0]    io_axiW_payload_strb,
  output              io_axiW_payload_last,
  input               io_axiB_valid,
  output              io_axiB_ready,
  input      [3:0]    io_axiB_payload_id,
  input      [1:0]    io_axiB_payload_resp,
  output              io_apDone,
  input               clk,
  input               reset
);
  reg                 buffer_1_io_push_valid;
  reg        [7:0]    buffer_1_io_push_payload;
  reg                 buffer_1_io_flush;
  wire                buffer_1_io_push_ready;
  wire                buffer_1_io_pop_valid;
  wire       [7:0]    buffer_1_io_pop_payload;
  wire       [5:0]    buffer_1_io_occupancy;
  wire       [5:0]    buffer_1_io_availability;
  wire       [8:0]    _zz_dataCounter_valueNext;
  wire       [0:0]    _zz_dataCounter_valueNext_1;
  wire       [8:0]    _zz_dataInCounter_valueNext;
  wire       [0:0]    _zz_dataInCounter_valueNext_1;
  wire       [7:0]    _zz_data255flag_valueNext;
  wire       [0:0]    _zz_data255flag_valueNext_1;
  wire       [31:0]   _zz_resdata;
  wire       [31:0]   _zz_regAwLen;
  wire       [39:0]   _zz_regAwAddr;
  wire       [31:0]   _zz_regAwAddr_1;
  wire       [31:0]   _zz_regAwLen_1;
  wire       [31:0]   _zz_when_AxiMasterWrite_l274;
  wire       [31:0]   _zz_when_AxiMasterWrite_l274_1;
  reg                 regApStart;
  reg        [31:0]   regWAO;
  reg        [31:0]   regALLWlen;
  reg                 dataCounter_willIncrement;
  reg                 dataCounter_willClear;
  reg        [8:0]    dataCounter_valueNext;
  reg        [8:0]    dataCounter_value;
  wire                dataCounter_willOverflowIfInc;
  wire                dataCounter_willOverflow;
  reg                 dataInCounter_willIncrement;
  reg                 dataInCounter_willClear;
  reg        [8:0]    dataInCounter_valueNext;
  reg        [8:0]    dataInCounter_value;
  wire                dataInCounter_willOverflowIfInc;
  wire                dataInCounter_willOverflow;
  reg                 data255flag_willIncrement;
  reg                 data255flag_willClear;
  reg        [7:0]    data255flag_valueNext;
  reg        [7:0]    data255flag_value;
  wire                data255flag_willOverflowIfInc;
  wire                data255flag_willOverflow;
  reg        [31:0]   regAwAddr;
  reg        [7:0]    regAwLen;
  reg                 regConfigFinish;
  reg                 regwlast;
  reg                 regApDone;
  wire       [31:0]   resdata;
  reg                 firstIn;
  reg                 regWriteFinish;
  wire                when_AxiMasterWrite_l186;
  wire                when_AxiMasterWrite_l197;
  wire                when_AxiMasterWrite_l198;
  wire                when_AxiMasterWrite_l209;
  wire                when_AxiMasterWrite_l218;
  wire                when_AxiMasterWrite_l256;
  wire                when_AxiMasterWrite_l274;
  wire                when_AxiMasterWrite_l276;

  assign _zz_dataCounter_valueNext_1 = dataCounter_willIncrement;
  assign _zz_dataCounter_valueNext = {8'd0, _zz_dataCounter_valueNext_1};
  assign _zz_dataInCounter_valueNext_1 = dataInCounter_willIncrement;
  assign _zz_dataInCounter_valueNext = {8'd0, _zz_dataInCounter_valueNext_1};
  assign _zz_data255flag_valueNext_1 = data255flag_willIncrement;
  assign _zz_data255flag_valueNext = {7'd0, _zz_data255flag_valueNext_1};
  assign _zz_resdata = {23'd0, dataCounter_value};
  assign _zz_regAwLen = (regWAO - 32'h00000001);
  assign _zz_regAwAddr = ({8'd0,_zz_regAwAddr_1} <<< 8);
  assign _zz_regAwAddr_1 = (regAwAddr + 32'h00000001);
  assign _zz_regAwLen_1 = (resdata - 32'h00000001);
  assign _zz_when_AxiMasterWrite_l274 = {23'd0, dataCounter_value};
  assign _zz_when_AxiMasterWrite_l274_1 = (io_Wlen - 32'h00000002);
  StreamFifo buffer_1 (
    .io_push_valid      (buffer_1_io_push_valid    ), //i
    .io_push_ready      (buffer_1_io_push_ready    ), //o
    .io_push_payload    (buffer_1_io_push_payload  ), //i
    .io_pop_valid       (buffer_1_io_pop_valid     ), //o
    .io_pop_ready       (io_axiW_ready             ), //i
    .io_pop_payload     (buffer_1_io_pop_payload   ), //o
    .io_flush           (buffer_1_io_flush         ), //i
    .io_occupancy       (buffer_1_io_occupancy     ), //o
    .io_availability    (buffer_1_io_availability  ), //o
    .clk                (clk                       ), //i
    .reset              (reset                     )  //i
  );
  always @(*) begin
    dataCounter_willIncrement = 1'b0;
    if(when_AxiMasterWrite_l256) begin
      dataCounter_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    dataCounter_willClear = 1'b0;
    if(dataCounter_willOverflow) begin
      dataCounter_willClear = 1'b1;
    end
  end

  assign dataCounter_willOverflowIfInc = (dataCounter_value == 9'h12b);
  assign dataCounter_willOverflow = (dataCounter_willOverflowIfInc && dataCounter_willIncrement);
  always @(*) begin
    if(dataCounter_willOverflow) begin
      dataCounter_valueNext = 9'h0;
    end else begin
      dataCounter_valueNext = (dataCounter_value + _zz_dataCounter_valueNext);
    end
    if(dataCounter_willClear) begin
      dataCounter_valueNext = 9'h0;
    end
  end

  always @(*) begin
    dataInCounter_willIncrement = 1'b0;
    if(when_AxiMasterWrite_l186) begin
      dataInCounter_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    dataInCounter_willClear = 1'b0;
    if(dataInCounter_willOverflow) begin
      dataInCounter_willClear = 1'b1;
    end
  end

  assign dataInCounter_willOverflowIfInc = (dataInCounter_value == 9'h12b);
  assign dataInCounter_willOverflow = (dataInCounter_willOverflowIfInc && dataInCounter_willIncrement);
  always @(*) begin
    if(dataInCounter_willOverflow) begin
      dataInCounter_valueNext = 9'h0;
    end else begin
      dataInCounter_valueNext = (dataInCounter_value + _zz_dataInCounter_valueNext);
    end
    if(dataInCounter_willClear) begin
      dataInCounter_valueNext = 9'h0;
    end
  end

  always @(*) begin
    data255flag_willIncrement = 1'b0;
    if(when_AxiMasterWrite_l256) begin
      data255flag_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    data255flag_willClear = 1'b0;
    if(dataCounter_willOverflow) begin
      data255flag_willClear = 1'b1;
    end
  end

  assign data255flag_willOverflowIfInc = (data255flag_value == 8'hff);
  assign data255flag_willOverflow = (data255flag_willOverflowIfInc && data255flag_willIncrement);
  always @(*) begin
    data255flag_valueNext = (data255flag_value + _zz_data255flag_valueNext);
    if(data255flag_willClear) begin
      data255flag_valueNext = 8'h0;
    end
  end

  assign io_data_in_ready = (((buffer_1_io_availability != 6'h0) && (! regWriteFinish)) && regApStart);
  assign when_AxiMasterWrite_l186 = (io_data_in_valid && io_data_in_ready);
  always @(*) begin
    if(when_AxiMasterWrite_l186) begin
      buffer_1_io_push_valid = 1'b1;
    end else begin
      buffer_1_io_push_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l186) begin
      buffer_1_io_push_payload = io_data_in_payload;
    end else begin
      buffer_1_io_push_payload = 8'h0;
    end
  end

  assign resdata = (regALLWlen - _zz_resdata);
  assign io_axiB_ready = 1'b1;
  assign when_AxiMasterWrite_l197 = (((regApStart && (! regConfigFinish)) && (! regWriteFinish)) && (firstIn || (io_axiB_valid && io_axiB_ready)));
  assign when_AxiMasterWrite_l198 = (regALLWlen < 32'h00000100);
  assign when_AxiMasterWrite_l209 = (resdata < 32'h00000100);
  assign when_AxiMasterWrite_l218 = ((regApStart && (! regApDone)) && regConfigFinish);
  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_valid = 1'b1;
    end else begin
      io_axiAW_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_addr = regAwAddr;
    end else begin
      io_axiAW_payload_addr = 32'h0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_burst = 2'b01;
    end else begin
      io_axiAW_payload_burst = 2'b00;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_size = 3'b000;
    end else begin
      io_axiAW_payload_size = 3'b000;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_len = regAwLen;
    end else begin
      io_axiAW_payload_len = 8'h0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_id = 4'b0000;
    end else begin
      io_axiAW_payload_id = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_lock = 1'b0;
    end else begin
      io_axiAW_payload_lock = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_region = 4'b0000;
    end else begin
      io_axiAW_payload_region = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_cache = 4'b0000;
    end else begin
      io_axiAW_payload_cache = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_qos = 4'b0000;
    end else begin
      io_axiAW_payload_qos = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_user = 1'b0;
    end else begin
      io_axiAW_payload_user = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterWrite_l218) begin
      io_axiAW_payload_prot = 3'b000;
    end else begin
      io_axiAW_payload_prot = 3'b000;
    end
  end

  assign io_axiW_valid = buffer_1_io_pop_valid;
  assign io_axiW_payload_data = buffer_1_io_pop_payload;
  assign io_axiW_payload_last = (regwlast && (io_axiW_valid && io_axiW_ready));
  assign io_axiW_payload_strb = 1'b1;
  assign io_apDone = regApDone;
  assign when_AxiMasterWrite_l256 = (io_axiW_valid && io_axiW_ready);
  always @(*) begin
    buffer_1_io_flush = 1'b0;
    if(regApDone) begin
      buffer_1_io_flush = 1'b1;
    end
  end

  assign when_AxiMasterWrite_l274 = (((dataCounter_value != 9'h0) && ((data255flag_value == 8'hfe) || (_zz_when_AxiMasterWrite_l274 == _zz_when_AxiMasterWrite_l274_1))) && (io_axiW_valid && io_axiW_ready));
  assign when_AxiMasterWrite_l276 = (regwlast && (io_axiW_valid && io_axiW_ready));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      regApStart <= 1'b0;
      regWAO <= 32'h0;
      regALLWlen <= 32'h0;
      dataCounter_value <= 9'h0;
      dataInCounter_value <= 9'h0;
      data255flag_value <= 8'h0;
      regAwAddr <= io_WAddrOffset;
      regAwLen <= 8'h0;
      regConfigFinish <= 1'b0;
      regwlast <= 1'b0;
      regApDone <= 1'b0;
      firstIn <= 1'b1;
      regWriteFinish <= 1'b0;
    end else begin
      regApStart <= io_apStart;
      regWAO <= io_WAddrOffset;
      regALLWlen <= io_Wlen;
      dataCounter_value <= dataCounter_valueNext;
      dataInCounter_value <= dataInCounter_valueNext;
      data255flag_value <= data255flag_valueNext;
      if(when_AxiMasterWrite_l197) begin
        if(when_AxiMasterWrite_l198) begin
          regAwAddr <= regWAO;
          regAwLen <= _zz_regAwLen[7:0];
          firstIn <= 1'b0;
        end else begin
          if(firstIn) begin
            regAwAddr <= regWAO;
            firstIn <= 1'b0;
          end else begin
            regAwAddr <= _zz_regAwAddr[31:0];
          end
          if(when_AxiMasterWrite_l209) begin
            regAwLen <= _zz_regAwLen_1[7:0];
          end else begin
            regAwLen <= 8'hff;
          end
        end
        regConfigFinish <= 1'b1;
      end
      if(data255flag_willOverflow) begin
        regConfigFinish <= 1'b0;
      end
      if(dataCounter_willOverflow) begin
        regApDone <= 1'b1;
      end
      if(dataInCounter_willOverflow) begin
        regWriteFinish <= 1'b1;
      end
      if(when_AxiMasterWrite_l274) begin
        regwlast <= 1'b1;
      end else begin
        if(when_AxiMasterWrite_l276) begin
          regwlast <= 1'b0;
        end
      end
      if(regApDone) begin
        regConfigFinish <= 1'b0;
        firstIn <= 1'b1;
        regApDone <= 1'b0;
        regWriteFinish <= 1'b0;
      end
    end
  end


endmodule

module AXI4MasterRead (
  output reg          io_dataOut_valid,
  input               io_dataOut_ready,
  output reg [7:0]    io_dataOut_payload,
  input               io_apStart,
  input      [31:0]   io_RAddrOffset,
  input      [31:0]   io_Rlen,
  output              io_apDone,
  output reg          io_axiAR_valid,
  input               io_axiAR_ready,
  output reg [31:0]   io_axiAR_payload_addr,
  output reg [3:0]    io_axiAR_payload_id,
  output reg [3:0]    io_axiAR_payload_region,
  output reg [7:0]    io_axiAR_payload_len,
  output reg [2:0]    io_axiAR_payload_size,
  output reg [1:0]    io_axiAR_payload_burst,
  output reg [0:0]    io_axiAR_payload_lock,
  output reg [3:0]    io_axiAR_payload_cache,
  output reg [3:0]    io_axiAR_payload_qos,
  output reg [0:0]    io_axiAR_payload_user,
  output reg [2:0]    io_axiAR_payload_prot,
  input               io_axiR_valid,
  output              io_axiR_ready,
  input      [7:0]    io_axiR_payload_data,
  input      [3:0]    io_axiR_payload_id,
  input      [1:0]    io_axiR_payload_resp,
  input               io_axiR_payload_last,
  input               clk,
  input               reset
);
  reg                 buffer_1_io_push_valid;
  reg        [7:0]    buffer_1_io_push_payload;
  reg                 buffer_1_io_pop_ready;
  wire                buffer_1_io_push_ready;
  wire                buffer_1_io_pop_valid;
  wire       [7:0]    buffer_1_io_pop_payload;
  wire       [5:0]    buffer_1_io_occupancy;
  wire       [5:0]    buffer_1_io_availability;
  wire       [8:0]    _zz_dataCounter_valueNext;
  wire       [0:0]    _zz_dataCounter_valueNext_1;
  wire       [31:0]   _zz_resdata;
  wire       [31:0]   _zz_regArLen;
  wire       [39:0]   _zz_regArAddr;
  wire       [31:0]   _zz_regArAddr_1;
  wire       [31:0]   _zz_regArLen_1;
  reg                 regApStart;
  reg        [31:0]   regRAO;
  reg        [31:0]   regALLRlen;
  reg                 dataCounter_willIncrement;
  wire                dataCounter_willClear;
  reg        [8:0]    dataCounter_valueNext;
  reg        [8:0]    dataCounter_value;
  wire                dataCounter_willOverflowIfInc;
  wire                dataCounter_willOverflow;
  reg        [31:0]   regArAddr;
  reg        [7:0]    regArLen;
  reg                 regConfigFinish;
  reg                 regApDone;
  reg                 firstIn;
  reg                 regReadFinsh;
  wire       [31:0]   resdata;
  wire                when_AxiMasterRead_l47;
  wire                when_AxiMasterRead_l48;
  wire                when_AxiMasterRead_l59;
  wire                when_AxiMasterRead_l67;
  wire                when_AxiMasterRead_l97;
  wire                when_AxiMasterRead_l108;
  wire                when_AxiMasterRead_l118;

  assign _zz_dataCounter_valueNext_1 = dataCounter_willIncrement;
  assign _zz_dataCounter_valueNext = {8'd0, _zz_dataCounter_valueNext_1};
  assign _zz_resdata = {23'd0, dataCounter_value};
  assign _zz_regArLen = (regRAO - 32'h00000001);
  assign _zz_regArAddr = ({8'd0,_zz_regArAddr_1} <<< 8);
  assign _zz_regArAddr_1 = (regArAddr + 32'h00000001);
  assign _zz_regArLen_1 = (resdata - 32'h00000001);
  StreamFifo buffer_1 (
    .io_push_valid      (buffer_1_io_push_valid    ), //i
    .io_push_ready      (buffer_1_io_push_ready    ), //o
    .io_push_payload    (buffer_1_io_push_payload  ), //i
    .io_pop_valid       (buffer_1_io_pop_valid     ), //o
    .io_pop_ready       (buffer_1_io_pop_ready     ), //i
    .io_pop_payload     (buffer_1_io_pop_payload   ), //o
    .io_flush           (1'b0                      ), //i
    .io_occupancy       (buffer_1_io_occupancy     ), //o
    .io_availability    (buffer_1_io_availability  ), //o
    .clk                (clk                       ), //i
    .reset              (reset                     )  //i
  );
  always @(*) begin
    dataCounter_willIncrement = 1'b0;
    if(when_AxiMasterRead_l97) begin
      dataCounter_willIncrement = 1'b1;
    end
  end

  assign dataCounter_willClear = 1'b0;
  assign dataCounter_willOverflowIfInc = (dataCounter_value == 9'h12b);
  assign dataCounter_willOverflow = (dataCounter_willOverflowIfInc && dataCounter_willIncrement);
  always @(*) begin
    if(dataCounter_willOverflow) begin
      dataCounter_valueNext = 9'h0;
    end else begin
      dataCounter_valueNext = (dataCounter_value + _zz_dataCounter_valueNext);
    end
    if(dataCounter_willClear) begin
      dataCounter_valueNext = 9'h0;
    end
  end

  assign resdata = (regALLRlen - _zz_resdata);
  assign when_AxiMasterRead_l47 = ((regApStart && (! regConfigFinish)) && (! regReadFinsh));
  assign when_AxiMasterRead_l48 = (regALLRlen < 32'h00000100);
  assign when_AxiMasterRead_l59 = (resdata < 32'h00000100);
  assign when_AxiMasterRead_l67 = ((regApStart && regConfigFinish) && (! regReadFinsh));
  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_valid = 1'b1;
    end else begin
      io_axiAR_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_addr = regArAddr;
    end else begin
      io_axiAR_payload_addr = 32'h0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_burst = 2'b01;
    end else begin
      io_axiAR_payload_burst = 2'b00;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_size = 3'b000;
    end else begin
      io_axiAR_payload_size = 3'b000;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_len = regArLen;
    end else begin
      io_axiAR_payload_len = 8'h0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_id = 4'b0000;
    end else begin
      io_axiAR_payload_id = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_lock = 1'b0;
    end else begin
      io_axiAR_payload_lock = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_region = 4'b0000;
    end else begin
      io_axiAR_payload_region = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_cache = 4'b0000;
    end else begin
      io_axiAR_payload_cache = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_qos = 4'b0000;
    end else begin
      io_axiAR_payload_qos = 4'b0000;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_user = 1'b0;
    end else begin
      io_axiAR_payload_user = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l67) begin
      io_axiAR_payload_prot = 3'b000;
    end else begin
      io_axiAR_payload_prot = 3'b000;
    end
  end

  assign io_axiR_ready = (buffer_1_io_availability != 6'h0);
  assign when_AxiMasterRead_l97 = (io_axiR_valid && io_axiR_ready);
  always @(*) begin
    if(when_AxiMasterRead_l97) begin
      buffer_1_io_push_valid = 1'b1;
    end else begin
      buffer_1_io_push_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l97) begin
      buffer_1_io_push_payload = io_axiR_payload_data;
    end else begin
      buffer_1_io_push_payload = 8'h0;
    end
  end

  assign when_AxiMasterRead_l108 = (buffer_1_io_occupancy != 6'h0);
  always @(*) begin
    if(when_AxiMasterRead_l108) begin
      io_dataOut_valid = buffer_1_io_pop_valid;
    end else begin
      io_dataOut_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l108) begin
      buffer_1_io_pop_ready = io_dataOut_ready;
    end else begin
      buffer_1_io_pop_ready = 1'b0;
    end
  end

  always @(*) begin
    if(when_AxiMasterRead_l108) begin
      io_dataOut_payload = buffer_1_io_pop_payload;
    end else begin
      io_dataOut_payload = 8'h0;
    end
  end

  assign when_AxiMasterRead_l118 = ((regReadFinsh && (buffer_1_io_occupancy == 6'h01)) && (io_dataOut_valid && io_dataOut_ready));
  assign io_apDone = regApDone;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      regApStart <= 1'b0;
      regRAO <= 32'h0;
      regALLRlen <= 32'h0;
      dataCounter_value <= 9'h0;
      regArAddr <= io_RAddrOffset;
      regArLen <= 8'h0;
      regConfigFinish <= 1'b0;
      regApDone <= 1'b0;
      firstIn <= 1'b1;
      regReadFinsh <= 1'b0;
    end else begin
      regApStart <= io_apStart;
      regRAO <= io_RAddrOffset;
      regALLRlen <= io_Rlen;
      dataCounter_value <= dataCounter_valueNext;
      if(when_AxiMasterRead_l47) begin
        if(when_AxiMasterRead_l48) begin
          regArAddr <= regRAO;
          regArLen <= _zz_regArLen[7:0];
          firstIn <= 1'b0;
        end else begin
          if(firstIn) begin
            regArAddr <= regRAO;
            firstIn <= 1'b0;
          end else begin
            regArAddr <= _zz_regArAddr[31:0];
          end
          if(when_AxiMasterRead_l59) begin
            regArLen <= _zz_regArLen_1[7:0];
          end else begin
            regArLen <= 8'hff;
          end
        end
        regConfigFinish <= 1'b1;
      end
      if(io_axiR_payload_last) begin
        regConfigFinish <= 1'b0;
      end
      if(dataCounter_willOverflow) begin
        regReadFinsh <= 1'b1;
      end
      if(when_AxiMasterRead_l118) begin
        regApDone <= 1'b1;
      end
      if(regApDone) begin
        regConfigFinish <= 1'b0;
        firstIn <= 1'b1;
        regReadFinsh <= 1'b0;
        regApDone <= 1'b0;
      end
    end
  end


endmodule

module Axi4_transmission (
  input               axiSignal_aw_valid,
  output              axiSignal_aw_ready,
  input      [31:0]   axiSignal_aw_payload_addr,
  input      [3:0]    axiSignal_aw_payload_id,
  input      [3:0]    axiSignal_aw_payload_region,
  input      [7:0]    axiSignal_aw_payload_len,
  input      [2:0]    axiSignal_aw_payload_size,
  input      [1:0]    axiSignal_aw_payload_burst,
  input      [0:0]    axiSignal_aw_payload_lock,
  input      [3:0]    axiSignal_aw_payload_cache,
  input      [3:0]    axiSignal_aw_payload_qos,
  input      [0:0]    axiSignal_aw_payload_user,
  input      [2:0]    axiSignal_aw_payload_prot,
  input               axiSignal_w_valid,
  output              axiSignal_w_ready,
  input      [7:0]    axiSignal_w_payload_data,
  input      [0:0]    axiSignal_w_payload_strb,
  input               axiSignal_w_payload_last,
  output              axiSignal_b_valid,
  input               axiSignal_b_ready,
  output     [3:0]    axiSignal_b_payload_id,
  output     [1:0]    axiSignal_b_payload_resp,
  input               axiSignal_ar_valid,
  output              axiSignal_ar_ready,
  input      [31:0]   axiSignal_ar_payload_addr,
  input      [3:0]    axiSignal_ar_payload_id,
  input      [3:0]    axiSignal_ar_payload_region,
  input      [7:0]    axiSignal_ar_payload_len,
  input      [2:0]    axiSignal_ar_payload_size,
  input      [1:0]    axiSignal_ar_payload_burst,
  input      [0:0]    axiSignal_ar_payload_lock,
  input      [3:0]    axiSignal_ar_payload_cache,
  input      [3:0]    axiSignal_ar_payload_qos,
  input      [0:0]    axiSignal_ar_payload_user,
  input      [2:0]    axiSignal_ar_payload_prot,
  output reg          axiSignal_r_valid,
  input               axiSignal_r_ready,
  output     [7:0]    axiSignal_r_payload_data,
  output     [3:0]    axiSignal_r_payload_id,
  output     [1:0]    axiSignal_r_payload_resp,
  output              axiSignal_r_payload_last,
  input               apstart,
  input               axireset,
  input               clk,
  input               reset
);
  wire       [12:0]   _zz_rFireCounter_valueNext;
  wire       [0:0]    _zz_rFireCounter_valueNext_1;
  wire       [31:0]   _zz_regAwAddr;
  wire       [11:0]   _zz__zz_1;
  reg        [7:0]    _zz__zz_regVec_0;
  wire       [11:0]   _zz__zz_regVec_0_1;
  reg        [7:0]    _zz__zz_regVec_0_1_1;
  wire       [11:0]   _zz_Axi4Incr_base;
  wire       [11:0]   _zz_Axi4Incr_base_1;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [31:0]   _zz_regArAddr;
  reg        [7:0]    _zz_axiSignal_r_payload_data;
  wire       [11:0]   _zz_axiSignal_r_payload_data_1;
  wire       [11:0]   _zz_Axi4Incr_base_1_1;
  wire       [11:0]   _zz_Axi4Incr_base_1_2;
  wire       [11:0]   _zz_Axi4Incr_baseIncr_1;
  reg        [11:0]   _zz_Axi4Incr_result_1;
  wire       [12:0]   _zz_when_Axi4_transmission_l177;
  wire       [12:0]   _zz_when_Axi4_transmission_l182;
  wire       [7:0]    _zz_when_Axi4_transmission_l182_1;
  reg        [7:0]    regVec_0;
  reg        [7:0]    regVec_1;
  reg        [7:0]    regVec_2;
  reg        [7:0]    regVec_3;
  reg        [7:0]    regVec_4;
  reg        [7:0]    regVec_5;
  reg        [7:0]    regVec_6;
  reg        [7:0]    regVec_7;
  reg        [7:0]    regVec_8;
  reg        [7:0]    regVec_9;
  reg        [7:0]    regVec_10;
  reg        [7:0]    regVec_11;
  reg        [7:0]    regVec_12;
  reg        [7:0]    regVec_13;
  reg        [7:0]    regVec_14;
  reg        [7:0]    regVec_15;
  reg        [7:0]    regVec_16;
  reg        [7:0]    regVec_17;
  reg        [7:0]    regVec_18;
  reg        [7:0]    regVec_19;
  reg        [7:0]    regVec_20;
  reg        [7:0]    regVec_21;
  reg        [7:0]    regVec_22;
  reg        [7:0]    regVec_23;
  reg        [7:0]    regVec_24;
  reg        [7:0]    regVec_25;
  reg        [7:0]    regVec_26;
  reg        [7:0]    regVec_27;
  reg        [7:0]    regVec_28;
  reg        [7:0]    regVec_29;
  reg        [7:0]    regVec_30;
  reg        [7:0]    regVec_31;
  reg        [7:0]    regVec_32;
  reg        [7:0]    regVec_33;
  reg        [7:0]    regVec_34;
  reg        [7:0]    regVec_35;
  reg        [7:0]    regVec_36;
  reg        [7:0]    regVec_37;
  reg        [7:0]    regVec_38;
  reg        [7:0]    regVec_39;
  reg        [7:0]    regVec_40;
  reg        [7:0]    regVec_41;
  reg        [7:0]    regVec_42;
  reg        [7:0]    regVec_43;
  reg        [7:0]    regVec_44;
  reg        [7:0]    regVec_45;
  reg        [7:0]    regVec_46;
  reg        [7:0]    regVec_47;
  reg        [7:0]    regVec_48;
  reg        [7:0]    regVec_49;
  reg        [7:0]    regVec_50;
  reg        [7:0]    regVec_51;
  reg        [7:0]    regVec_52;
  reg        [7:0]    regVec_53;
  reg        [7:0]    regVec_54;
  reg        [7:0]    regVec_55;
  reg        [7:0]    regVec_56;
  reg        [7:0]    regVec_57;
  reg        [7:0]    regVec_58;
  reg        [7:0]    regVec_59;
  reg        [7:0]    regVec_60;
  reg        [7:0]    regVec_61;
  reg        [7:0]    regVec_62;
  reg        [7:0]    regVec_63;
  reg        [7:0]    regVec_64;
  reg        [7:0]    regVec_65;
  reg        [7:0]    regVec_66;
  reg        [7:0]    regVec_67;
  reg        [7:0]    regVec_68;
  reg        [7:0]    regVec_69;
  reg        [7:0]    regVec_70;
  reg        [7:0]    regVec_71;
  reg        [7:0]    regVec_72;
  reg        [7:0]    regVec_73;
  reg        [7:0]    regVec_74;
  reg        [7:0]    regVec_75;
  reg        [7:0]    regVec_76;
  reg        [7:0]    regVec_77;
  reg        [7:0]    regVec_78;
  reg        [7:0]    regVec_79;
  reg        [7:0]    regVec_80;
  reg        [7:0]    regVec_81;
  reg        [7:0]    regVec_82;
  reg        [7:0]    regVec_83;
  reg        [7:0]    regVec_84;
  reg        [7:0]    regVec_85;
  reg        [7:0]    regVec_86;
  reg        [7:0]    regVec_87;
  reg        [7:0]    regVec_88;
  reg        [7:0]    regVec_89;
  reg        [7:0]    regVec_90;
  reg        [7:0]    regVec_91;
  reg        [7:0]    regVec_92;
  reg        [7:0]    regVec_93;
  reg        [7:0]    regVec_94;
  reg        [7:0]    regVec_95;
  reg        [7:0]    regVec_96;
  reg        [7:0]    regVec_97;
  reg        [7:0]    regVec_98;
  reg        [7:0]    regVec_99;
  reg        [7:0]    regVec_100;
  reg        [7:0]    regVec_101;
  reg        [7:0]    regVec_102;
  reg        [7:0]    regVec_103;
  reg        [7:0]    regVec_104;
  reg        [7:0]    regVec_105;
  reg        [7:0]    regVec_106;
  reg        [7:0]    regVec_107;
  reg        [7:0]    regVec_108;
  reg        [7:0]    regVec_109;
  reg        [7:0]    regVec_110;
  reg        [7:0]    regVec_111;
  reg        [7:0]    regVec_112;
  reg        [7:0]    regVec_113;
  reg        [7:0]    regVec_114;
  reg        [7:0]    regVec_115;
  reg        [7:0]    regVec_116;
  reg        [7:0]    regVec_117;
  reg        [7:0]    regVec_118;
  reg        [7:0]    regVec_119;
  reg        [7:0]    regVec_120;
  reg        [7:0]    regVec_121;
  reg        [7:0]    regVec_122;
  reg        [7:0]    regVec_123;
  reg        [7:0]    regVec_124;
  reg        [7:0]    regVec_125;
  reg        [7:0]    regVec_126;
  reg        [7:0]    regVec_127;
  reg        [7:0]    regVec_128;
  reg        [7:0]    regVec_129;
  reg        [7:0]    regVec_130;
  reg        [7:0]    regVec_131;
  reg        [7:0]    regVec_132;
  reg        [7:0]    regVec_133;
  reg        [7:0]    regVec_134;
  reg        [7:0]    regVec_135;
  reg        [7:0]    regVec_136;
  reg        [7:0]    regVec_137;
  reg        [7:0]    regVec_138;
  reg        [7:0]    regVec_139;
  reg        [7:0]    regVec_140;
  reg        [7:0]    regVec_141;
  reg        [7:0]    regVec_142;
  reg        [7:0]    regVec_143;
  reg        [7:0]    regVec_144;
  reg        [7:0]    regVec_145;
  reg        [7:0]    regVec_146;
  reg        [7:0]    regVec_147;
  reg        [7:0]    regVec_148;
  reg        [7:0]    regVec_149;
  reg        [7:0]    regVec_150;
  reg        [7:0]    regVec_151;
  reg        [7:0]    regVec_152;
  reg        [7:0]    regVec_153;
  reg        [7:0]    regVec_154;
  reg        [7:0]    regVec_155;
  reg        [7:0]    regVec_156;
  reg        [7:0]    regVec_157;
  reg        [7:0]    regVec_158;
  reg        [7:0]    regVec_159;
  reg        [7:0]    regVec_160;
  reg        [7:0]    regVec_161;
  reg        [7:0]    regVec_162;
  reg        [7:0]    regVec_163;
  reg        [7:0]    regVec_164;
  reg        [7:0]    regVec_165;
  reg        [7:0]    regVec_166;
  reg        [7:0]    regVec_167;
  reg        [7:0]    regVec_168;
  reg        [7:0]    regVec_169;
  reg        [7:0]    regVec_170;
  reg        [7:0]    regVec_171;
  reg        [7:0]    regVec_172;
  reg        [7:0]    regVec_173;
  reg        [7:0]    regVec_174;
  reg        [7:0]    regVec_175;
  reg        [7:0]    regVec_176;
  reg        [7:0]    regVec_177;
  reg        [7:0]    regVec_178;
  reg        [7:0]    regVec_179;
  reg        [7:0]    regVec_180;
  reg        [7:0]    regVec_181;
  reg        [7:0]    regVec_182;
  reg        [7:0]    regVec_183;
  reg        [7:0]    regVec_184;
  reg        [7:0]    regVec_185;
  reg        [7:0]    regVec_186;
  reg        [7:0]    regVec_187;
  reg        [7:0]    regVec_188;
  reg        [7:0]    regVec_189;
  reg        [7:0]    regVec_190;
  reg        [7:0]    regVec_191;
  reg        [7:0]    regVec_192;
  reg        [7:0]    regVec_193;
  reg        [7:0]    regVec_194;
  reg        [7:0]    regVec_195;
  reg        [7:0]    regVec_196;
  reg        [7:0]    regVec_197;
  reg        [7:0]    regVec_198;
  reg        [7:0]    regVec_199;
  reg        [7:0]    regVec_200;
  reg        [7:0]    regVec_201;
  reg        [7:0]    regVec_202;
  reg        [7:0]    regVec_203;
  reg        [7:0]    regVec_204;
  reg        [7:0]    regVec_205;
  reg        [7:0]    regVec_206;
  reg        [7:0]    regVec_207;
  reg        [7:0]    regVec_208;
  reg        [7:0]    regVec_209;
  reg        [7:0]    regVec_210;
  reg        [7:0]    regVec_211;
  reg        [7:0]    regVec_212;
  reg        [7:0]    regVec_213;
  reg        [7:0]    regVec_214;
  reg        [7:0]    regVec_215;
  reg        [7:0]    regVec_216;
  reg        [7:0]    regVec_217;
  reg        [7:0]    regVec_218;
  reg        [7:0]    regVec_219;
  reg        [7:0]    regVec_220;
  reg        [7:0]    regVec_221;
  reg        [7:0]    regVec_222;
  reg        [7:0]    regVec_223;
  reg        [7:0]    regVec_224;
  reg        [7:0]    regVec_225;
  reg        [7:0]    regVec_226;
  reg        [7:0]    regVec_227;
  reg        [7:0]    regVec_228;
  reg        [7:0]    regVec_229;
  reg        [7:0]    regVec_230;
  reg        [7:0]    regVec_231;
  reg        [7:0]    regVec_232;
  reg        [7:0]    regVec_233;
  reg        [7:0]    regVec_234;
  reg        [7:0]    regVec_235;
  reg        [7:0]    regVec_236;
  reg        [7:0]    regVec_237;
  reg        [7:0]    regVec_238;
  reg        [7:0]    regVec_239;
  reg        [7:0]    regVec_240;
  reg        [7:0]    regVec_241;
  reg        [7:0]    regVec_242;
  reg        [7:0]    regVec_243;
  reg        [7:0]    regVec_244;
  reg        [7:0]    regVec_245;
  reg        [7:0]    regVec_246;
  reg        [7:0]    regVec_247;
  reg        [7:0]    regVec_248;
  reg        [7:0]    regVec_249;
  reg        [7:0]    regVec_250;
  reg        [7:0]    regVec_251;
  reg        [7:0]    regVec_252;
  reg        [7:0]    regVec_253;
  reg        [7:0]    regVec_254;
  reg        [7:0]    regVec_255;
  reg        [7:0]    regVec_256;
  reg        [7:0]    regVec_257;
  reg        [7:0]    regVec_258;
  reg        [7:0]    regVec_259;
  reg        [7:0]    regVec_260;
  reg        [7:0]    regVec_261;
  reg        [7:0]    regVec_262;
  reg        [7:0]    regVec_263;
  reg        [7:0]    regVec_264;
  reg        [7:0]    regVec_265;
  reg        [7:0]    regVec_266;
  reg        [7:0]    regVec_267;
  reg        [7:0]    regVec_268;
  reg        [7:0]    regVec_269;
  reg        [7:0]    regVec_270;
  reg        [7:0]    regVec_271;
  reg        [7:0]    regVec_272;
  reg        [7:0]    regVec_273;
  reg        [7:0]    regVec_274;
  reg        [7:0]    regVec_275;
  reg        [7:0]    regVec_276;
  reg        [7:0]    regVec_277;
  reg        [7:0]    regVec_278;
  reg        [7:0]    regVec_279;
  reg        [7:0]    regVec_280;
  reg        [7:0]    regVec_281;
  reg        [7:0]    regVec_282;
  reg        [7:0]    regVec_283;
  reg        [7:0]    regVec_284;
  reg        [7:0]    regVec_285;
  reg        [7:0]    regVec_286;
  reg        [7:0]    regVec_287;
  reg        [7:0]    regVec_288;
  reg        [7:0]    regVec_289;
  reg        [7:0]    regVec_290;
  reg        [7:0]    regVec_291;
  reg        [7:0]    regVec_292;
  reg        [7:0]    regVec_293;
  reg        [7:0]    regVec_294;
  reg        [7:0]    regVec_295;
  reg        [7:0]    regVec_296;
  reg        [7:0]    regVec_297;
  reg        [7:0]    regVec_298;
  reg        [7:0]    regVec_299;
  reg        [7:0]    regVec_300;
  reg        [7:0]    regVec_301;
  reg        [7:0]    regVec_302;
  reg        [7:0]    regVec_303;
  reg        [7:0]    regVec_304;
  reg        [7:0]    regVec_305;
  reg        [7:0]    regVec_306;
  reg        [7:0]    regVec_307;
  reg        [7:0]    regVec_308;
  reg        [7:0]    regVec_309;
  reg        [7:0]    regVec_310;
  reg        [7:0]    regVec_311;
  reg        [7:0]    regVec_312;
  reg        [7:0]    regVec_313;
  reg        [7:0]    regVec_314;
  reg        [7:0]    regVec_315;
  reg        [7:0]    regVec_316;
  reg        [7:0]    regVec_317;
  reg        [7:0]    regVec_318;
  reg        [7:0]    regVec_319;
  reg        [7:0]    regVec_320;
  reg        [7:0]    regVec_321;
  reg        [7:0]    regVec_322;
  reg        [7:0]    regVec_323;
  reg        [7:0]    regVec_324;
  reg        [7:0]    regVec_325;
  reg        [7:0]    regVec_326;
  reg        [7:0]    regVec_327;
  reg        [7:0]    regVec_328;
  reg        [7:0]    regVec_329;
  reg        [7:0]    regVec_330;
  reg        [7:0]    regVec_331;
  reg        [7:0]    regVec_332;
  reg        [7:0]    regVec_333;
  reg        [7:0]    regVec_334;
  reg        [7:0]    regVec_335;
  reg        [7:0]    regVec_336;
  reg        [7:0]    regVec_337;
  reg        [7:0]    regVec_338;
  reg        [7:0]    regVec_339;
  reg        [7:0]    regVec_340;
  reg        [7:0]    regVec_341;
  reg        [7:0]    regVec_342;
  reg        [7:0]    regVec_343;
  reg        [7:0]    regVec_344;
  reg        [7:0]    regVec_345;
  reg        [7:0]    regVec_346;
  reg        [7:0]    regVec_347;
  reg        [7:0]    regVec_348;
  reg        [7:0]    regVec_349;
  reg        [7:0]    regVec_350;
  reg        [7:0]    regVec_351;
  reg        [7:0]    regVec_352;
  reg        [7:0]    regVec_353;
  reg        [7:0]    regVec_354;
  reg        [7:0]    regVec_355;
  reg        [7:0]    regVec_356;
  reg        [7:0]    regVec_357;
  reg        [7:0]    regVec_358;
  reg        [7:0]    regVec_359;
  reg        [7:0]    regVec_360;
  reg        [7:0]    regVec_361;
  reg        [7:0]    regVec_362;
  reg        [7:0]    regVec_363;
  reg        [7:0]    regVec_364;
  reg        [7:0]    regVec_365;
  reg        [7:0]    regVec_366;
  reg        [7:0]    regVec_367;
  reg        [7:0]    regVec_368;
  reg        [7:0]    regVec_369;
  reg        [7:0]    regVec_370;
  reg        [7:0]    regVec_371;
  reg        [7:0]    regVec_372;
  reg        [7:0]    regVec_373;
  reg        [7:0]    regVec_374;
  reg        [7:0]    regVec_375;
  reg        [7:0]    regVec_376;
  reg        [7:0]    regVec_377;
  reg        [7:0]    regVec_378;
  reg        [7:0]    regVec_379;
  reg        [7:0]    regVec_380;
  reg        [7:0]    regVec_381;
  reg        [7:0]    regVec_382;
  reg        [7:0]    regVec_383;
  reg        [7:0]    regVec_384;
  reg        [7:0]    regVec_385;
  reg        [7:0]    regVec_386;
  reg        [7:0]    regVec_387;
  reg        [7:0]    regVec_388;
  reg        [7:0]    regVec_389;
  reg        [7:0]    regVec_390;
  reg        [7:0]    regVec_391;
  reg        [7:0]    regVec_392;
  reg        [7:0]    regVec_393;
  reg        [7:0]    regVec_394;
  reg        [7:0]    regVec_395;
  reg        [7:0]    regVec_396;
  reg        [7:0]    regVec_397;
  reg        [7:0]    regVec_398;
  reg        [7:0]    regVec_399;
  reg        [7:0]    regVec_400;
  reg        [7:0]    regVec_401;
  reg        [7:0]    regVec_402;
  reg        [7:0]    regVec_403;
  reg        [7:0]    regVec_404;
  reg        [7:0]    regVec_405;
  reg        [7:0]    regVec_406;
  reg        [7:0]    regVec_407;
  reg        [7:0]    regVec_408;
  reg        [7:0]    regVec_409;
  reg        [7:0]    regVec_410;
  reg        [7:0]    regVec_411;
  reg        [7:0]    regVec_412;
  reg        [7:0]    regVec_413;
  reg        [7:0]    regVec_414;
  reg        [7:0]    regVec_415;
  reg        [7:0]    regVec_416;
  reg        [7:0]    regVec_417;
  reg        [7:0]    regVec_418;
  reg        [7:0]    regVec_419;
  reg        [7:0]    regVec_420;
  reg        [7:0]    regVec_421;
  reg        [7:0]    regVec_422;
  reg        [7:0]    regVec_423;
  reg        [7:0]    regVec_424;
  reg        [7:0]    regVec_425;
  reg        [7:0]    regVec_426;
  reg        [7:0]    regVec_427;
  reg        [7:0]    regVec_428;
  reg        [7:0]    regVec_429;
  reg        [7:0]    regVec_430;
  reg        [7:0]    regVec_431;
  reg        [7:0]    regVec_432;
  reg        [7:0]    regVec_433;
  reg        [7:0]    regVec_434;
  reg        [7:0]    regVec_435;
  reg        [7:0]    regVec_436;
  reg        [7:0]    regVec_437;
  reg        [7:0]    regVec_438;
  reg        [7:0]    regVec_439;
  reg        [7:0]    regVec_440;
  reg        [7:0]    regVec_441;
  reg        [7:0]    regVec_442;
  reg        [7:0]    regVec_443;
  reg        [7:0]    regVec_444;
  reg        [7:0]    regVec_445;
  reg        [7:0]    regVec_446;
  reg        [7:0]    regVec_447;
  reg        [7:0]    regVec_448;
  reg        [7:0]    regVec_449;
  reg        [7:0]    regVec_450;
  reg        [7:0]    regVec_451;
  reg        [7:0]    regVec_452;
  reg        [7:0]    regVec_453;
  reg        [7:0]    regVec_454;
  reg        [7:0]    regVec_455;
  reg        [7:0]    regVec_456;
  reg        [7:0]    regVec_457;
  reg        [7:0]    regVec_458;
  reg        [7:0]    regVec_459;
  reg        [7:0]    regVec_460;
  reg        [7:0]    regVec_461;
  reg        [7:0]    regVec_462;
  reg        [7:0]    regVec_463;
  reg        [7:0]    regVec_464;
  reg        [7:0]    regVec_465;
  reg        [7:0]    regVec_466;
  reg        [7:0]    regVec_467;
  reg        [7:0]    regVec_468;
  reg        [7:0]    regVec_469;
  reg        [7:0]    regVec_470;
  reg        [7:0]    regVec_471;
  reg        [7:0]    regVec_472;
  reg        [7:0]    regVec_473;
  reg        [7:0]    regVec_474;
  reg        [7:0]    regVec_475;
  reg        [7:0]    regVec_476;
  reg        [7:0]    regVec_477;
  reg        [7:0]    regVec_478;
  reg        [7:0]    regVec_479;
  reg        [7:0]    regVec_480;
  reg        [7:0]    regVec_481;
  reg        [7:0]    regVec_482;
  reg        [7:0]    regVec_483;
  reg        [7:0]    regVec_484;
  reg        [7:0]    regVec_485;
  reg        [7:0]    regVec_486;
  reg        [7:0]    regVec_487;
  reg        [7:0]    regVec_488;
  reg        [7:0]    regVec_489;
  reg        [7:0]    regVec_490;
  reg        [7:0]    regVec_491;
  reg        [7:0]    regVec_492;
  reg        [7:0]    regVec_493;
  reg        [7:0]    regVec_494;
  reg        [7:0]    regVec_495;
  reg        [7:0]    regVec_496;
  reg        [7:0]    regVec_497;
  reg        [7:0]    regVec_498;
  reg        [7:0]    regVec_499;
  reg        [7:0]    regVec_500;
  reg        [7:0]    regVec_501;
  reg        [7:0]    regVec_502;
  reg        [7:0]    regVec_503;
  reg        [7:0]    regVec_504;
  reg        [7:0]    regVec_505;
  reg        [7:0]    regVec_506;
  reg        [7:0]    regVec_507;
  reg        [7:0]    regVec_508;
  reg        [7:0]    regVec_509;
  reg        [7:0]    regVec_510;
  reg        [7:0]    regVec_511;
  reg        [7:0]    regVec_512;
  reg        [7:0]    regVec_513;
  reg        [7:0]    regVec_514;
  reg        [7:0]    regVec_515;
  reg        [7:0]    regVec_516;
  reg        [7:0]    regVec_517;
  reg        [7:0]    regVec_518;
  reg        [7:0]    regVec_519;
  reg        [7:0]    regVec_520;
  reg        [7:0]    regVec_521;
  reg        [7:0]    regVec_522;
  reg        [7:0]    regVec_523;
  reg        [7:0]    regVec_524;
  reg        [7:0]    regVec_525;
  reg        [7:0]    regVec_526;
  reg        [7:0]    regVec_527;
  reg        [7:0]    regVec_528;
  reg        [7:0]    regVec_529;
  reg        [7:0]    regVec_530;
  reg        [7:0]    regVec_531;
  reg        [7:0]    regVec_532;
  reg        [7:0]    regVec_533;
  reg        [7:0]    regVec_534;
  reg        [7:0]    regVec_535;
  reg        [7:0]    regVec_536;
  reg        [7:0]    regVec_537;
  reg        [7:0]    regVec_538;
  reg        [7:0]    regVec_539;
  reg        [7:0]    regVec_540;
  reg        [7:0]    regVec_541;
  reg        [7:0]    regVec_542;
  reg        [7:0]    regVec_543;
  reg        [7:0]    regVec_544;
  reg        [7:0]    regVec_545;
  reg        [7:0]    regVec_546;
  reg        [7:0]    regVec_547;
  reg        [7:0]    regVec_548;
  reg        [7:0]    regVec_549;
  reg        [7:0]    regVec_550;
  reg        [7:0]    regVec_551;
  reg        [7:0]    regVec_552;
  reg        [7:0]    regVec_553;
  reg        [7:0]    regVec_554;
  reg        [7:0]    regVec_555;
  reg        [7:0]    regVec_556;
  reg        [7:0]    regVec_557;
  reg        [7:0]    regVec_558;
  reg        [7:0]    regVec_559;
  reg        [7:0]    regVec_560;
  reg        [7:0]    regVec_561;
  reg        [7:0]    regVec_562;
  reg        [7:0]    regVec_563;
  reg        [7:0]    regVec_564;
  reg        [7:0]    regVec_565;
  reg        [7:0]    regVec_566;
  reg        [7:0]    regVec_567;
  reg        [7:0]    regVec_568;
  reg        [7:0]    regVec_569;
  reg        [7:0]    regVec_570;
  reg        [7:0]    regVec_571;
  reg        [7:0]    regVec_572;
  reg        [7:0]    regVec_573;
  reg        [7:0]    regVec_574;
  reg        [7:0]    regVec_575;
  reg        [7:0]    regVec_576;
  reg        [7:0]    regVec_577;
  reg        [7:0]    regVec_578;
  reg        [7:0]    regVec_579;
  reg        [7:0]    regVec_580;
  reg        [7:0]    regVec_581;
  reg        [7:0]    regVec_582;
  reg        [7:0]    regVec_583;
  reg        [7:0]    regVec_584;
  reg        [7:0]    regVec_585;
  reg        [7:0]    regVec_586;
  reg        [7:0]    regVec_587;
  reg        [7:0]    regVec_588;
  reg        [7:0]    regVec_589;
  reg        [7:0]    regVec_590;
  reg        [7:0]    regVec_591;
  reg        [7:0]    regVec_592;
  reg        [7:0]    regVec_593;
  reg        [7:0]    regVec_594;
  reg        [7:0]    regVec_595;
  reg        [7:0]    regVec_596;
  reg        [7:0]    regVec_597;
  reg        [7:0]    regVec_598;
  reg        [7:0]    regVec_599;
  reg        [7:0]    regVec_600;
  reg        [7:0]    regVec_601;
  reg        [7:0]    regVec_602;
  reg        [7:0]    regVec_603;
  reg        [7:0]    regVec_604;
  reg        [7:0]    regVec_605;
  reg        [7:0]    regVec_606;
  reg        [7:0]    regVec_607;
  reg        [7:0]    regVec_608;
  reg        [7:0]    regVec_609;
  reg        [7:0]    regVec_610;
  reg        [7:0]    regVec_611;
  reg        [7:0]    regVec_612;
  reg        [7:0]    regVec_613;
  reg        [7:0]    regVec_614;
  reg        [7:0]    regVec_615;
  reg        [7:0]    regVec_616;
  reg        [7:0]    regVec_617;
  reg        [7:0]    regVec_618;
  reg        [7:0]    regVec_619;
  reg        [7:0]    regVec_620;
  reg        [7:0]    regVec_621;
  reg        [7:0]    regVec_622;
  reg        [7:0]    regVec_623;
  reg        [7:0]    regVec_624;
  reg        [7:0]    regVec_625;
  reg        [7:0]    regVec_626;
  reg        [7:0]    regVec_627;
  reg        [7:0]    regVec_628;
  reg        [7:0]    regVec_629;
  reg        [7:0]    regVec_630;
  reg        [7:0]    regVec_631;
  reg        [7:0]    regVec_632;
  reg        [7:0]    regVec_633;
  reg        [7:0]    regVec_634;
  reg        [7:0]    regVec_635;
  reg        [7:0]    regVec_636;
  reg        [7:0]    regVec_637;
  reg        [7:0]    regVec_638;
  reg        [7:0]    regVec_639;
  reg        [7:0]    regVec_640;
  reg        [7:0]    regVec_641;
  reg        [7:0]    regVec_642;
  reg        [7:0]    regVec_643;
  reg        [7:0]    regVec_644;
  reg        [7:0]    regVec_645;
  reg        [7:0]    regVec_646;
  reg        [7:0]    regVec_647;
  reg        [7:0]    regVec_648;
  reg        [7:0]    regVec_649;
  reg        [7:0]    regVec_650;
  reg        [7:0]    regVec_651;
  reg        [7:0]    regVec_652;
  reg        [7:0]    regVec_653;
  reg        [7:0]    regVec_654;
  reg        [7:0]    regVec_655;
  reg        [7:0]    regVec_656;
  reg        [7:0]    regVec_657;
  reg        [7:0]    regVec_658;
  reg        [7:0]    regVec_659;
  reg        [7:0]    regVec_660;
  reg        [7:0]    regVec_661;
  reg        [7:0]    regVec_662;
  reg        [7:0]    regVec_663;
  reg        [7:0]    regVec_664;
  reg        [7:0]    regVec_665;
  reg        [7:0]    regVec_666;
  reg        [7:0]    regVec_667;
  reg        [7:0]    regVec_668;
  reg        [7:0]    regVec_669;
  reg        [7:0]    regVec_670;
  reg        [7:0]    regVec_671;
  reg        [7:0]    regVec_672;
  reg        [7:0]    regVec_673;
  reg        [7:0]    regVec_674;
  reg        [7:0]    regVec_675;
  reg        [7:0]    regVec_676;
  reg        [7:0]    regVec_677;
  reg        [7:0]    regVec_678;
  reg        [7:0]    regVec_679;
  reg        [7:0]    regVec_680;
  reg        [7:0]    regVec_681;
  reg        [7:0]    regVec_682;
  reg        [7:0]    regVec_683;
  reg        [7:0]    regVec_684;
  reg        [7:0]    regVec_685;
  reg        [7:0]    regVec_686;
  reg        [7:0]    regVec_687;
  reg        [7:0]    regVec_688;
  reg        [7:0]    regVec_689;
  reg        [7:0]    regVec_690;
  reg        [7:0]    regVec_691;
  reg        [7:0]    regVec_692;
  reg        [7:0]    regVec_693;
  reg        [7:0]    regVec_694;
  reg        [7:0]    regVec_695;
  reg        [7:0]    regVec_696;
  reg        [7:0]    regVec_697;
  reg        [7:0]    regVec_698;
  reg        [7:0]    regVec_699;
  reg        [7:0]    regVec_700;
  reg        [7:0]    regVec_701;
  reg        [7:0]    regVec_702;
  reg        [7:0]    regVec_703;
  reg        [7:0]    regVec_704;
  reg        [7:0]    regVec_705;
  reg        [7:0]    regVec_706;
  reg        [7:0]    regVec_707;
  reg        [7:0]    regVec_708;
  reg        [7:0]    regVec_709;
  reg        [7:0]    regVec_710;
  reg        [7:0]    regVec_711;
  reg        [7:0]    regVec_712;
  reg        [7:0]    regVec_713;
  reg        [7:0]    regVec_714;
  reg        [7:0]    regVec_715;
  reg        [7:0]    regVec_716;
  reg        [7:0]    regVec_717;
  reg        [7:0]    regVec_718;
  reg        [7:0]    regVec_719;
  reg        [7:0]    regVec_720;
  reg        [7:0]    regVec_721;
  reg        [7:0]    regVec_722;
  reg        [7:0]    regVec_723;
  reg        [7:0]    regVec_724;
  reg        [7:0]    regVec_725;
  reg        [7:0]    regVec_726;
  reg        [7:0]    regVec_727;
  reg        [7:0]    regVec_728;
  reg        [7:0]    regVec_729;
  reg        [7:0]    regVec_730;
  reg        [7:0]    regVec_731;
  reg        [7:0]    regVec_732;
  reg        [7:0]    regVec_733;
  reg        [7:0]    regVec_734;
  reg        [7:0]    regVec_735;
  reg        [7:0]    regVec_736;
  reg        [7:0]    regVec_737;
  reg        [7:0]    regVec_738;
  reg        [7:0]    regVec_739;
  reg        [7:0]    regVec_740;
  reg        [7:0]    regVec_741;
  reg        [7:0]    regVec_742;
  reg        [7:0]    regVec_743;
  reg        [7:0]    regVec_744;
  reg        [7:0]    regVec_745;
  reg        [7:0]    regVec_746;
  reg        [7:0]    regVec_747;
  reg        [7:0]    regVec_748;
  reg        [7:0]    regVec_749;
  reg        [7:0]    regVec_750;
  reg        [7:0]    regVec_751;
  reg        [7:0]    regVec_752;
  reg        [7:0]    regVec_753;
  reg        [7:0]    regVec_754;
  reg        [7:0]    regVec_755;
  reg        [7:0]    regVec_756;
  reg        [7:0]    regVec_757;
  reg        [7:0]    regVec_758;
  reg        [7:0]    regVec_759;
  reg        [7:0]    regVec_760;
  reg        [7:0]    regVec_761;
  reg        [7:0]    regVec_762;
  reg        [7:0]    regVec_763;
  reg        [7:0]    regVec_764;
  reg        [7:0]    regVec_765;
  reg        [7:0]    regVec_766;
  reg        [7:0]    regVec_767;
  reg        [7:0]    regVec_768;
  reg        [7:0]    regVec_769;
  reg        [7:0]    regVec_770;
  reg        [7:0]    regVec_771;
  reg        [7:0]    regVec_772;
  reg        [7:0]    regVec_773;
  reg        [7:0]    regVec_774;
  reg        [7:0]    regVec_775;
  reg        [7:0]    regVec_776;
  reg        [7:0]    regVec_777;
  reg        [7:0]    regVec_778;
  reg        [7:0]    regVec_779;
  reg        [7:0]    regVec_780;
  reg        [7:0]    regVec_781;
  reg        [7:0]    regVec_782;
  reg        [7:0]    regVec_783;
  reg        [7:0]    regVec_784;
  reg        [7:0]    regVec_785;
  reg        [7:0]    regVec_786;
  reg        [7:0]    regVec_787;
  reg        [7:0]    regVec_788;
  reg        [7:0]    regVec_789;
  reg        [7:0]    regVec_790;
  reg        [7:0]    regVec_791;
  reg        [7:0]    regVec_792;
  reg        [7:0]    regVec_793;
  reg        [7:0]    regVec_794;
  reg        [7:0]    regVec_795;
  reg        [7:0]    regVec_796;
  reg        [7:0]    regVec_797;
  reg        [7:0]    regVec_798;
  reg        [7:0]    regVec_799;
  reg        [7:0]    regVec_800;
  reg        [7:0]    regVec_801;
  reg        [7:0]    regVec_802;
  reg        [7:0]    regVec_803;
  reg        [7:0]    regVec_804;
  reg        [7:0]    regVec_805;
  reg        [7:0]    regVec_806;
  reg        [7:0]    regVec_807;
  reg        [7:0]    regVec_808;
  reg        [7:0]    regVec_809;
  reg        [7:0]    regVec_810;
  reg        [7:0]    regVec_811;
  reg        [7:0]    regVec_812;
  reg        [7:0]    regVec_813;
  reg        [7:0]    regVec_814;
  reg        [7:0]    regVec_815;
  reg        [7:0]    regVec_816;
  reg        [7:0]    regVec_817;
  reg        [7:0]    regVec_818;
  reg        [7:0]    regVec_819;
  reg        [7:0]    regVec_820;
  reg        [7:0]    regVec_821;
  reg        [7:0]    regVec_822;
  reg        [7:0]    regVec_823;
  reg        [7:0]    regVec_824;
  reg        [7:0]    regVec_825;
  reg        [7:0]    regVec_826;
  reg        [7:0]    regVec_827;
  reg        [7:0]    regVec_828;
  reg        [7:0]    regVec_829;
  reg        [7:0]    regVec_830;
  reg        [7:0]    regVec_831;
  reg        [7:0]    regVec_832;
  reg        [7:0]    regVec_833;
  reg        [7:0]    regVec_834;
  reg        [7:0]    regVec_835;
  reg        [7:0]    regVec_836;
  reg        [7:0]    regVec_837;
  reg        [7:0]    regVec_838;
  reg        [7:0]    regVec_839;
  reg        [7:0]    regVec_840;
  reg        [7:0]    regVec_841;
  reg        [7:0]    regVec_842;
  reg        [7:0]    regVec_843;
  reg        [7:0]    regVec_844;
  reg        [7:0]    regVec_845;
  reg        [7:0]    regVec_846;
  reg        [7:0]    regVec_847;
  reg        [7:0]    regVec_848;
  reg        [7:0]    regVec_849;
  reg        [7:0]    regVec_850;
  reg        [7:0]    regVec_851;
  reg        [7:0]    regVec_852;
  reg        [7:0]    regVec_853;
  reg        [7:0]    regVec_854;
  reg        [7:0]    regVec_855;
  reg        [7:0]    regVec_856;
  reg        [7:0]    regVec_857;
  reg        [7:0]    regVec_858;
  reg        [7:0]    regVec_859;
  reg        [7:0]    regVec_860;
  reg        [7:0]    regVec_861;
  reg        [7:0]    regVec_862;
  reg        [7:0]    regVec_863;
  reg        [7:0]    regVec_864;
  reg        [7:0]    regVec_865;
  reg        [7:0]    regVec_866;
  reg        [7:0]    regVec_867;
  reg        [7:0]    regVec_868;
  reg        [7:0]    regVec_869;
  reg        [7:0]    regVec_870;
  reg        [7:0]    regVec_871;
  reg        [7:0]    regVec_872;
  reg        [7:0]    regVec_873;
  reg        [7:0]    regVec_874;
  reg        [7:0]    regVec_875;
  reg        [7:0]    regVec_876;
  reg        [7:0]    regVec_877;
  reg        [7:0]    regVec_878;
  reg        [7:0]    regVec_879;
  reg        [7:0]    regVec_880;
  reg        [7:0]    regVec_881;
  reg        [7:0]    regVec_882;
  reg        [7:0]    regVec_883;
  reg        [7:0]    regVec_884;
  reg        [7:0]    regVec_885;
  reg        [7:0]    regVec_886;
  reg        [7:0]    regVec_887;
  reg        [7:0]    regVec_888;
  reg        [7:0]    regVec_889;
  reg        [7:0]    regVec_890;
  reg        [7:0]    regVec_891;
  reg        [7:0]    regVec_892;
  reg        [7:0]    regVec_893;
  reg        [7:0]    regVec_894;
  reg        [7:0]    regVec_895;
  reg        [7:0]    regVec_896;
  reg        [7:0]    regVec_897;
  reg        [7:0]    regVec_898;
  reg        [7:0]    regVec_899;
  reg        [7:0]    regVec_900;
  reg        [7:0]    regVec_901;
  reg        [7:0]    regVec_902;
  reg        [7:0]    regVec_903;
  reg        [7:0]    regVec_904;
  reg        [7:0]    regVec_905;
  reg        [7:0]    regVec_906;
  reg        [7:0]    regVec_907;
  reg        [7:0]    regVec_908;
  reg        [7:0]    regVec_909;
  reg        [7:0]    regVec_910;
  reg        [7:0]    regVec_911;
  reg        [7:0]    regVec_912;
  reg        [7:0]    regVec_913;
  reg        [7:0]    regVec_914;
  reg        [7:0]    regVec_915;
  reg        [7:0]    regVec_916;
  reg        [7:0]    regVec_917;
  reg        [7:0]    regVec_918;
  reg        [7:0]    regVec_919;
  reg        [7:0]    regVec_920;
  reg        [7:0]    regVec_921;
  reg        [7:0]    regVec_922;
  reg        [7:0]    regVec_923;
  reg        [7:0]    regVec_924;
  reg        [7:0]    regVec_925;
  reg        [7:0]    regVec_926;
  reg        [7:0]    regVec_927;
  reg        [7:0]    regVec_928;
  reg        [7:0]    regVec_929;
  reg        [7:0]    regVec_930;
  reg        [7:0]    regVec_931;
  reg        [7:0]    regVec_932;
  reg        [7:0]    regVec_933;
  reg        [7:0]    regVec_934;
  reg        [7:0]    regVec_935;
  reg        [7:0]    regVec_936;
  reg        [7:0]    regVec_937;
  reg        [7:0]    regVec_938;
  reg        [7:0]    regVec_939;
  reg        [7:0]    regVec_940;
  reg        [7:0]    regVec_941;
  reg        [7:0]    regVec_942;
  reg        [7:0]    regVec_943;
  reg        [7:0]    regVec_944;
  reg        [7:0]    regVec_945;
  reg        [7:0]    regVec_946;
  reg        [7:0]    regVec_947;
  reg        [7:0]    regVec_948;
  reg        [7:0]    regVec_949;
  reg        [7:0]    regVec_950;
  reg        [7:0]    regVec_951;
  reg        [7:0]    regVec_952;
  reg        [7:0]    regVec_953;
  reg        [7:0]    regVec_954;
  reg        [7:0]    regVec_955;
  reg        [7:0]    regVec_956;
  reg        [7:0]    regVec_957;
  reg        [7:0]    regVec_958;
  reg        [7:0]    regVec_959;
  reg        [7:0]    regVec_960;
  reg        [7:0]    regVec_961;
  reg        [7:0]    regVec_962;
  reg        [7:0]    regVec_963;
  reg        [7:0]    regVec_964;
  reg        [7:0]    regVec_965;
  reg        [7:0]    regVec_966;
  reg        [7:0]    regVec_967;
  reg        [7:0]    regVec_968;
  reg        [7:0]    regVec_969;
  reg        [7:0]    regVec_970;
  reg        [7:0]    regVec_971;
  reg        [7:0]    regVec_972;
  reg        [7:0]    regVec_973;
  reg        [7:0]    regVec_974;
  reg        [7:0]    regVec_975;
  reg        [7:0]    regVec_976;
  reg        [7:0]    regVec_977;
  reg        [7:0]    regVec_978;
  reg        [7:0]    regVec_979;
  reg        [7:0]    regVec_980;
  reg        [7:0]    regVec_981;
  reg        [7:0]    regVec_982;
  reg        [7:0]    regVec_983;
  reg        [7:0]    regVec_984;
  reg        [7:0]    regVec_985;
  reg        [7:0]    regVec_986;
  reg        [7:0]    regVec_987;
  reg        [7:0]    regVec_988;
  reg        [7:0]    regVec_989;
  reg        [7:0]    regVec_990;
  reg        [7:0]    regVec_991;
  reg        [7:0]    regVec_992;
  reg        [7:0]    regVec_993;
  reg        [7:0]    regVec_994;
  reg        [7:0]    regVec_995;
  reg        [7:0]    regVec_996;
  reg        [7:0]    regVec_997;
  reg        [7:0]    regVec_998;
  reg        [7:0]    regVec_999;
  reg        [7:0]    regVec_1000;
  reg        [7:0]    regVec_1001;
  reg        [7:0]    regVec_1002;
  reg        [7:0]    regVec_1003;
  reg        [7:0]    regVec_1004;
  reg        [7:0]    regVec_1005;
  reg        [7:0]    regVec_1006;
  reg        [7:0]    regVec_1007;
  reg        [7:0]    regVec_1008;
  reg        [7:0]    regVec_1009;
  reg        [7:0]    regVec_1010;
  reg        [7:0]    regVec_1011;
  reg        [7:0]    regVec_1012;
  reg        [7:0]    regVec_1013;
  reg        [7:0]    regVec_1014;
  reg        [7:0]    regVec_1015;
  reg        [7:0]    regVec_1016;
  reg        [7:0]    regVec_1017;
  reg        [7:0]    regVec_1018;
  reg        [7:0]    regVec_1019;
  reg        [7:0]    regVec_1020;
  reg        [7:0]    regVec_1021;
  reg        [7:0]    regVec_1022;
  reg        [7:0]    regVec_1023;
  reg        [7:0]    regVec_1024;
  reg        [7:0]    regVec_1025;
  reg        [7:0]    regVec_1026;
  reg        [7:0]    regVec_1027;
  reg        [7:0]    regVec_1028;
  reg        [7:0]    regVec_1029;
  reg        [7:0]    regVec_1030;
  reg        [7:0]    regVec_1031;
  reg        [7:0]    regVec_1032;
  reg        [7:0]    regVec_1033;
  reg        [7:0]    regVec_1034;
  reg        [7:0]    regVec_1035;
  reg        [7:0]    regVec_1036;
  reg        [7:0]    regVec_1037;
  reg        [7:0]    regVec_1038;
  reg        [7:0]    regVec_1039;
  reg        [7:0]    regVec_1040;
  reg        [7:0]    regVec_1041;
  reg        [7:0]    regVec_1042;
  reg        [7:0]    regVec_1043;
  reg        [7:0]    regVec_1044;
  reg        [7:0]    regVec_1045;
  reg        [7:0]    regVec_1046;
  reg        [7:0]    regVec_1047;
  reg        [7:0]    regVec_1048;
  reg        [7:0]    regVec_1049;
  reg        [7:0]    regVec_1050;
  reg        [7:0]    regVec_1051;
  reg        [7:0]    regVec_1052;
  reg        [7:0]    regVec_1053;
  reg        [7:0]    regVec_1054;
  reg        [7:0]    regVec_1055;
  reg        [7:0]    regVec_1056;
  reg        [7:0]    regVec_1057;
  reg        [7:0]    regVec_1058;
  reg        [7:0]    regVec_1059;
  reg        [7:0]    regVec_1060;
  reg        [7:0]    regVec_1061;
  reg        [7:0]    regVec_1062;
  reg        [7:0]    regVec_1063;
  reg        [7:0]    regVec_1064;
  reg        [7:0]    regVec_1065;
  reg        [7:0]    regVec_1066;
  reg        [7:0]    regVec_1067;
  reg        [7:0]    regVec_1068;
  reg        [7:0]    regVec_1069;
  reg        [7:0]    regVec_1070;
  reg        [7:0]    regVec_1071;
  reg        [7:0]    regVec_1072;
  reg        [7:0]    regVec_1073;
  reg        [7:0]    regVec_1074;
  reg        [7:0]    regVec_1075;
  reg        [7:0]    regVec_1076;
  reg        [7:0]    regVec_1077;
  reg        [7:0]    regVec_1078;
  reg        [7:0]    regVec_1079;
  reg        [7:0]    regVec_1080;
  reg        [7:0]    regVec_1081;
  reg        [7:0]    regVec_1082;
  reg        [7:0]    regVec_1083;
  reg        [7:0]    regVec_1084;
  reg        [7:0]    regVec_1085;
  reg        [7:0]    regVec_1086;
  reg        [7:0]    regVec_1087;
  reg        [7:0]    regVec_1088;
  reg        [7:0]    regVec_1089;
  reg        [7:0]    regVec_1090;
  reg        [7:0]    regVec_1091;
  reg        [7:0]    regVec_1092;
  reg        [7:0]    regVec_1093;
  reg        [7:0]    regVec_1094;
  reg        [7:0]    regVec_1095;
  reg        [7:0]    regVec_1096;
  reg        [7:0]    regVec_1097;
  reg        [7:0]    regVec_1098;
  reg        [7:0]    regVec_1099;
  reg        [7:0]    regVec_1100;
  reg        [7:0]    regVec_1101;
  reg        [7:0]    regVec_1102;
  reg        [7:0]    regVec_1103;
  reg        [7:0]    regVec_1104;
  reg        [7:0]    regVec_1105;
  reg        [7:0]    regVec_1106;
  reg        [7:0]    regVec_1107;
  reg        [7:0]    regVec_1108;
  reg        [7:0]    regVec_1109;
  reg        [7:0]    regVec_1110;
  reg        [7:0]    regVec_1111;
  reg        [7:0]    regVec_1112;
  reg        [7:0]    regVec_1113;
  reg        [7:0]    regVec_1114;
  reg        [7:0]    regVec_1115;
  reg        [7:0]    regVec_1116;
  reg        [7:0]    regVec_1117;
  reg        [7:0]    regVec_1118;
  reg        [7:0]    regVec_1119;
  reg        [7:0]    regVec_1120;
  reg        [7:0]    regVec_1121;
  reg        [7:0]    regVec_1122;
  reg        [7:0]    regVec_1123;
  reg        [7:0]    regVec_1124;
  reg        [7:0]    regVec_1125;
  reg        [7:0]    regVec_1126;
  reg        [7:0]    regVec_1127;
  reg        [7:0]    regVec_1128;
  reg        [7:0]    regVec_1129;
  reg        [7:0]    regVec_1130;
  reg        [7:0]    regVec_1131;
  reg        [7:0]    regVec_1132;
  reg        [7:0]    regVec_1133;
  reg        [7:0]    regVec_1134;
  reg        [7:0]    regVec_1135;
  reg        [7:0]    regVec_1136;
  reg        [7:0]    regVec_1137;
  reg        [7:0]    regVec_1138;
  reg        [7:0]    regVec_1139;
  reg        [7:0]    regVec_1140;
  reg        [7:0]    regVec_1141;
  reg        [7:0]    regVec_1142;
  reg        [7:0]    regVec_1143;
  reg        [7:0]    regVec_1144;
  reg        [7:0]    regVec_1145;
  reg        [7:0]    regVec_1146;
  reg        [7:0]    regVec_1147;
  reg        [7:0]    regVec_1148;
  reg        [7:0]    regVec_1149;
  reg        [7:0]    regVec_1150;
  reg        [7:0]    regVec_1151;
  reg        [7:0]    regVec_1152;
  reg        [7:0]    regVec_1153;
  reg        [7:0]    regVec_1154;
  reg        [7:0]    regVec_1155;
  reg        [7:0]    regVec_1156;
  reg        [7:0]    regVec_1157;
  reg        [7:0]    regVec_1158;
  reg        [7:0]    regVec_1159;
  reg        [7:0]    regVec_1160;
  reg        [7:0]    regVec_1161;
  reg        [7:0]    regVec_1162;
  reg        [7:0]    regVec_1163;
  reg        [7:0]    regVec_1164;
  reg        [7:0]    regVec_1165;
  reg        [7:0]    regVec_1166;
  reg        [7:0]    regVec_1167;
  reg        [7:0]    regVec_1168;
  reg        [7:0]    regVec_1169;
  reg        [7:0]    regVec_1170;
  reg        [7:0]    regVec_1171;
  reg        [7:0]    regVec_1172;
  reg        [7:0]    regVec_1173;
  reg        [7:0]    regVec_1174;
  reg        [7:0]    regVec_1175;
  reg        [7:0]    regVec_1176;
  reg        [7:0]    regVec_1177;
  reg        [7:0]    regVec_1178;
  reg        [7:0]    regVec_1179;
  reg        [7:0]    regVec_1180;
  reg        [7:0]    regVec_1181;
  reg        [7:0]    regVec_1182;
  reg        [7:0]    regVec_1183;
  reg        [7:0]    regVec_1184;
  reg        [7:0]    regVec_1185;
  reg        [7:0]    regVec_1186;
  reg        [7:0]    regVec_1187;
  reg        [7:0]    regVec_1188;
  reg        [7:0]    regVec_1189;
  reg        [7:0]    regVec_1190;
  reg        [7:0]    regVec_1191;
  reg        [7:0]    regVec_1192;
  reg        [7:0]    regVec_1193;
  reg        [7:0]    regVec_1194;
  reg        [7:0]    regVec_1195;
  reg        [7:0]    regVec_1196;
  reg        [7:0]    regVec_1197;
  reg        [7:0]    regVec_1198;
  reg        [7:0]    regVec_1199;
  reg        [7:0]    regVec_1200;
  reg        [7:0]    regVec_1201;
  reg        [7:0]    regVec_1202;
  reg        [7:0]    regVec_1203;
  reg        [7:0]    regVec_1204;
  reg        [7:0]    regVec_1205;
  reg        [7:0]    regVec_1206;
  reg        [7:0]    regVec_1207;
  reg        [7:0]    regVec_1208;
  reg        [7:0]    regVec_1209;
  reg        [7:0]    regVec_1210;
  reg        [7:0]    regVec_1211;
  reg        [7:0]    regVec_1212;
  reg        [7:0]    regVec_1213;
  reg        [7:0]    regVec_1214;
  reg        [7:0]    regVec_1215;
  reg        [7:0]    regVec_1216;
  reg        [7:0]    regVec_1217;
  reg        [7:0]    regVec_1218;
  reg        [7:0]    regVec_1219;
  reg        [7:0]    regVec_1220;
  reg        [7:0]    regVec_1221;
  reg        [7:0]    regVec_1222;
  reg        [7:0]    regVec_1223;
  reg        [7:0]    regVec_1224;
  reg        [7:0]    regVec_1225;
  reg        [7:0]    regVec_1226;
  reg        [7:0]    regVec_1227;
  reg        [7:0]    regVec_1228;
  reg        [7:0]    regVec_1229;
  reg        [7:0]    regVec_1230;
  reg        [7:0]    regVec_1231;
  reg        [7:0]    regVec_1232;
  reg        [7:0]    regVec_1233;
  reg        [7:0]    regVec_1234;
  reg        [7:0]    regVec_1235;
  reg        [7:0]    regVec_1236;
  reg        [7:0]    regVec_1237;
  reg        [7:0]    regVec_1238;
  reg        [7:0]    regVec_1239;
  reg        [7:0]    regVec_1240;
  reg        [7:0]    regVec_1241;
  reg        [7:0]    regVec_1242;
  reg        [7:0]    regVec_1243;
  reg        [7:0]    regVec_1244;
  reg        [7:0]    regVec_1245;
  reg        [7:0]    regVec_1246;
  reg        [7:0]    regVec_1247;
  reg        [7:0]    regVec_1248;
  reg        [7:0]    regVec_1249;
  reg        [7:0]    regVec_1250;
  reg        [7:0]    regVec_1251;
  reg        [7:0]    regVec_1252;
  reg        [7:0]    regVec_1253;
  reg        [7:0]    regVec_1254;
  reg        [7:0]    regVec_1255;
  reg        [7:0]    regVec_1256;
  reg        [7:0]    regVec_1257;
  reg        [7:0]    regVec_1258;
  reg        [7:0]    regVec_1259;
  reg        [7:0]    regVec_1260;
  reg        [7:0]    regVec_1261;
  reg        [7:0]    regVec_1262;
  reg        [7:0]    regVec_1263;
  reg        [7:0]    regVec_1264;
  reg        [7:0]    regVec_1265;
  reg        [7:0]    regVec_1266;
  reg        [7:0]    regVec_1267;
  reg        [7:0]    regVec_1268;
  reg        [7:0]    regVec_1269;
  reg        [7:0]    regVec_1270;
  reg        [7:0]    regVec_1271;
  reg        [7:0]    regVec_1272;
  reg        [7:0]    regVec_1273;
  reg        [7:0]    regVec_1274;
  reg        [7:0]    regVec_1275;
  reg        [7:0]    regVec_1276;
  reg        [7:0]    regVec_1277;
  reg        [7:0]    regVec_1278;
  reg        [7:0]    regVec_1279;
  reg        [7:0]    regVec_1280;
  reg        [7:0]    regVec_1281;
  reg        [7:0]    regVec_1282;
  reg        [7:0]    regVec_1283;
  reg        [7:0]    regVec_1284;
  reg        [7:0]    regVec_1285;
  reg        [7:0]    regVec_1286;
  reg        [7:0]    regVec_1287;
  reg        [7:0]    regVec_1288;
  reg        [7:0]    regVec_1289;
  reg        [7:0]    regVec_1290;
  reg        [7:0]    regVec_1291;
  reg        [7:0]    regVec_1292;
  reg        [7:0]    regVec_1293;
  reg        [7:0]    regVec_1294;
  reg        [7:0]    regVec_1295;
  reg        [7:0]    regVec_1296;
  reg        [7:0]    regVec_1297;
  reg        [7:0]    regVec_1298;
  reg        [7:0]    regVec_1299;
  reg        [7:0]    regVec_1300;
  reg        [7:0]    regVec_1301;
  reg        [7:0]    regVec_1302;
  reg        [7:0]    regVec_1303;
  reg        [7:0]    regVec_1304;
  reg        [7:0]    regVec_1305;
  reg        [7:0]    regVec_1306;
  reg        [7:0]    regVec_1307;
  reg        [7:0]    regVec_1308;
  reg        [7:0]    regVec_1309;
  reg        [7:0]    regVec_1310;
  reg        [7:0]    regVec_1311;
  reg        [7:0]    regVec_1312;
  reg        [7:0]    regVec_1313;
  reg        [7:0]    regVec_1314;
  reg        [7:0]    regVec_1315;
  reg        [7:0]    regVec_1316;
  reg        [7:0]    regVec_1317;
  reg        [7:0]    regVec_1318;
  reg        [7:0]    regVec_1319;
  reg        [7:0]    regVec_1320;
  reg        [7:0]    regVec_1321;
  reg        [7:0]    regVec_1322;
  reg        [7:0]    regVec_1323;
  reg        [7:0]    regVec_1324;
  reg        [7:0]    regVec_1325;
  reg        [7:0]    regVec_1326;
  reg        [7:0]    regVec_1327;
  reg        [7:0]    regVec_1328;
  reg        [7:0]    regVec_1329;
  reg        [7:0]    regVec_1330;
  reg        [7:0]    regVec_1331;
  reg        [7:0]    regVec_1332;
  reg        [7:0]    regVec_1333;
  reg        [7:0]    regVec_1334;
  reg        [7:0]    regVec_1335;
  reg        [7:0]    regVec_1336;
  reg        [7:0]    regVec_1337;
  reg        [7:0]    regVec_1338;
  reg        [7:0]    regVec_1339;
  reg        [7:0]    regVec_1340;
  reg        [7:0]    regVec_1341;
  reg        [7:0]    regVec_1342;
  reg        [7:0]    regVec_1343;
  reg        [7:0]    regVec_1344;
  reg        [7:0]    regVec_1345;
  reg        [7:0]    regVec_1346;
  reg        [7:0]    regVec_1347;
  reg        [7:0]    regVec_1348;
  reg        [7:0]    regVec_1349;
  reg        [7:0]    regVec_1350;
  reg        [7:0]    regVec_1351;
  reg        [7:0]    regVec_1352;
  reg        [7:0]    regVec_1353;
  reg        [7:0]    regVec_1354;
  reg        [7:0]    regVec_1355;
  reg        [7:0]    regVec_1356;
  reg        [7:0]    regVec_1357;
  reg        [7:0]    regVec_1358;
  reg        [7:0]    regVec_1359;
  reg        [7:0]    regVec_1360;
  reg        [7:0]    regVec_1361;
  reg        [7:0]    regVec_1362;
  reg        [7:0]    regVec_1363;
  reg        [7:0]    regVec_1364;
  reg        [7:0]    regVec_1365;
  reg        [7:0]    regVec_1366;
  reg        [7:0]    regVec_1367;
  reg        [7:0]    regVec_1368;
  reg        [7:0]    regVec_1369;
  reg        [7:0]    regVec_1370;
  reg        [7:0]    regVec_1371;
  reg        [7:0]    regVec_1372;
  reg        [7:0]    regVec_1373;
  reg        [7:0]    regVec_1374;
  reg        [7:0]    regVec_1375;
  reg        [7:0]    regVec_1376;
  reg        [7:0]    regVec_1377;
  reg        [7:0]    regVec_1378;
  reg        [7:0]    regVec_1379;
  reg        [7:0]    regVec_1380;
  reg        [7:0]    regVec_1381;
  reg        [7:0]    regVec_1382;
  reg        [7:0]    regVec_1383;
  reg        [7:0]    regVec_1384;
  reg        [7:0]    regVec_1385;
  reg        [7:0]    regVec_1386;
  reg        [7:0]    regVec_1387;
  reg        [7:0]    regVec_1388;
  reg        [7:0]    regVec_1389;
  reg        [7:0]    regVec_1390;
  reg        [7:0]    regVec_1391;
  reg        [7:0]    regVec_1392;
  reg        [7:0]    regVec_1393;
  reg        [7:0]    regVec_1394;
  reg        [7:0]    regVec_1395;
  reg        [7:0]    regVec_1396;
  reg        [7:0]    regVec_1397;
  reg        [7:0]    regVec_1398;
  reg        [7:0]    regVec_1399;
  reg        [7:0]    regVec_1400;
  reg        [7:0]    regVec_1401;
  reg        [7:0]    regVec_1402;
  reg        [7:0]    regVec_1403;
  reg        [7:0]    regVec_1404;
  reg        [7:0]    regVec_1405;
  reg        [7:0]    regVec_1406;
  reg        [7:0]    regVec_1407;
  reg        [7:0]    regVec_1408;
  reg        [7:0]    regVec_1409;
  reg        [7:0]    regVec_1410;
  reg        [7:0]    regVec_1411;
  reg        [7:0]    regVec_1412;
  reg        [7:0]    regVec_1413;
  reg        [7:0]    regVec_1414;
  reg        [7:0]    regVec_1415;
  reg        [7:0]    regVec_1416;
  reg        [7:0]    regVec_1417;
  reg        [7:0]    regVec_1418;
  reg        [7:0]    regVec_1419;
  reg        [7:0]    regVec_1420;
  reg        [7:0]    regVec_1421;
  reg        [7:0]    regVec_1422;
  reg        [7:0]    regVec_1423;
  reg        [7:0]    regVec_1424;
  reg        [7:0]    regVec_1425;
  reg        [7:0]    regVec_1426;
  reg        [7:0]    regVec_1427;
  reg        [7:0]    regVec_1428;
  reg        [7:0]    regVec_1429;
  reg        [7:0]    regVec_1430;
  reg        [7:0]    regVec_1431;
  reg        [7:0]    regVec_1432;
  reg        [7:0]    regVec_1433;
  reg        [7:0]    regVec_1434;
  reg        [7:0]    regVec_1435;
  reg        [7:0]    regVec_1436;
  reg        [7:0]    regVec_1437;
  reg        [7:0]    regVec_1438;
  reg        [7:0]    regVec_1439;
  reg        [7:0]    regVec_1440;
  reg        [7:0]    regVec_1441;
  reg        [7:0]    regVec_1442;
  reg        [7:0]    regVec_1443;
  reg        [7:0]    regVec_1444;
  reg        [7:0]    regVec_1445;
  reg        [7:0]    regVec_1446;
  reg        [7:0]    regVec_1447;
  reg        [7:0]    regVec_1448;
  reg        [7:0]    regVec_1449;
  reg        [7:0]    regVec_1450;
  reg        [7:0]    regVec_1451;
  reg        [7:0]    regVec_1452;
  reg        [7:0]    regVec_1453;
  reg        [7:0]    regVec_1454;
  reg        [7:0]    regVec_1455;
  reg        [7:0]    regVec_1456;
  reg        [7:0]    regVec_1457;
  reg        [7:0]    regVec_1458;
  reg        [7:0]    regVec_1459;
  reg        [7:0]    regVec_1460;
  reg        [7:0]    regVec_1461;
  reg        [7:0]    regVec_1462;
  reg        [7:0]    regVec_1463;
  reg        [7:0]    regVec_1464;
  reg        [7:0]    regVec_1465;
  reg        [7:0]    regVec_1466;
  reg        [7:0]    regVec_1467;
  reg        [7:0]    regVec_1468;
  reg        [7:0]    regVec_1469;
  reg        [7:0]    regVec_1470;
  reg        [7:0]    regVec_1471;
  reg        [7:0]    regVec_1472;
  reg        [7:0]    regVec_1473;
  reg        [7:0]    regVec_1474;
  reg        [7:0]    regVec_1475;
  reg        [7:0]    regVec_1476;
  reg        [7:0]    regVec_1477;
  reg        [7:0]    regVec_1478;
  reg        [7:0]    regVec_1479;
  reg        [7:0]    regVec_1480;
  reg        [7:0]    regVec_1481;
  reg        [7:0]    regVec_1482;
  reg        [7:0]    regVec_1483;
  reg        [7:0]    regVec_1484;
  reg        [7:0]    regVec_1485;
  reg        [7:0]    regVec_1486;
  reg        [7:0]    regVec_1487;
  reg        [7:0]    regVec_1488;
  reg        [7:0]    regVec_1489;
  reg        [7:0]    regVec_1490;
  reg        [7:0]    regVec_1491;
  reg        [7:0]    regVec_1492;
  reg        [7:0]    regVec_1493;
  reg        [7:0]    regVec_1494;
  reg        [7:0]    regVec_1495;
  reg        [7:0]    regVec_1496;
  reg        [7:0]    regVec_1497;
  reg        [7:0]    regVec_1498;
  reg        [7:0]    regVec_1499;
  reg        [7:0]    regVec_1500;
  reg        [7:0]    regVec_1501;
  reg        [7:0]    regVec_1502;
  reg        [7:0]    regVec_1503;
  reg        [7:0]    regVec_1504;
  reg        [7:0]    regVec_1505;
  reg        [7:0]    regVec_1506;
  reg        [7:0]    regVec_1507;
  reg        [7:0]    regVec_1508;
  reg        [7:0]    regVec_1509;
  reg        [7:0]    regVec_1510;
  reg        [7:0]    regVec_1511;
  reg        [7:0]    regVec_1512;
  reg        [7:0]    regVec_1513;
  reg        [7:0]    regVec_1514;
  reg        [7:0]    regVec_1515;
  reg        [7:0]    regVec_1516;
  reg        [7:0]    regVec_1517;
  reg        [7:0]    regVec_1518;
  reg        [7:0]    regVec_1519;
  reg        [7:0]    regVec_1520;
  reg        [7:0]    regVec_1521;
  reg        [7:0]    regVec_1522;
  reg        [7:0]    regVec_1523;
  reg        [7:0]    regVec_1524;
  reg        [7:0]    regVec_1525;
  reg        [7:0]    regVec_1526;
  reg        [7:0]    regVec_1527;
  reg        [7:0]    regVec_1528;
  reg        [7:0]    regVec_1529;
  reg        [7:0]    regVec_1530;
  reg        [7:0]    regVec_1531;
  reg        [7:0]    regVec_1532;
  reg        [7:0]    regVec_1533;
  reg        [7:0]    regVec_1534;
  reg        [7:0]    regVec_1535;
  reg        [7:0]    regVec_1536;
  reg        [7:0]    regVec_1537;
  reg        [7:0]    regVec_1538;
  reg        [7:0]    regVec_1539;
  reg        [7:0]    regVec_1540;
  reg        [7:0]    regVec_1541;
  reg        [7:0]    regVec_1542;
  reg        [7:0]    regVec_1543;
  reg        [7:0]    regVec_1544;
  reg        [7:0]    regVec_1545;
  reg        [7:0]    regVec_1546;
  reg        [7:0]    regVec_1547;
  reg        [7:0]    regVec_1548;
  reg        [7:0]    regVec_1549;
  reg        [7:0]    regVec_1550;
  reg        [7:0]    regVec_1551;
  reg        [7:0]    regVec_1552;
  reg        [7:0]    regVec_1553;
  reg        [7:0]    regVec_1554;
  reg        [7:0]    regVec_1555;
  reg        [7:0]    regVec_1556;
  reg        [7:0]    regVec_1557;
  reg        [7:0]    regVec_1558;
  reg        [7:0]    regVec_1559;
  reg        [7:0]    regVec_1560;
  reg        [7:0]    regVec_1561;
  reg        [7:0]    regVec_1562;
  reg        [7:0]    regVec_1563;
  reg        [7:0]    regVec_1564;
  reg        [7:0]    regVec_1565;
  reg        [7:0]    regVec_1566;
  reg        [7:0]    regVec_1567;
  reg        [7:0]    regVec_1568;
  reg        [7:0]    regVec_1569;
  reg        [7:0]    regVec_1570;
  reg        [7:0]    regVec_1571;
  reg        [7:0]    regVec_1572;
  reg        [7:0]    regVec_1573;
  reg        [7:0]    regVec_1574;
  reg        [7:0]    regVec_1575;
  reg        [7:0]    regVec_1576;
  reg        [7:0]    regVec_1577;
  reg        [7:0]    regVec_1578;
  reg        [7:0]    regVec_1579;
  reg        [7:0]    regVec_1580;
  reg        [7:0]    regVec_1581;
  reg        [7:0]    regVec_1582;
  reg        [7:0]    regVec_1583;
  reg        [7:0]    regVec_1584;
  reg        [7:0]    regVec_1585;
  reg        [7:0]    regVec_1586;
  reg        [7:0]    regVec_1587;
  reg        [7:0]    regVec_1588;
  reg        [7:0]    regVec_1589;
  reg        [7:0]    regVec_1590;
  reg        [7:0]    regVec_1591;
  reg        [7:0]    regVec_1592;
  reg        [7:0]    regVec_1593;
  reg        [7:0]    regVec_1594;
  reg        [7:0]    regVec_1595;
  reg        [7:0]    regVec_1596;
  reg        [7:0]    regVec_1597;
  reg        [7:0]    regVec_1598;
  reg        [7:0]    regVec_1599;
  reg        [7:0]    regVec_1600;
  reg        [7:0]    regVec_1601;
  reg        [7:0]    regVec_1602;
  reg        [7:0]    regVec_1603;
  reg        [7:0]    regVec_1604;
  reg        [7:0]    regVec_1605;
  reg        [7:0]    regVec_1606;
  reg        [7:0]    regVec_1607;
  reg        [7:0]    regVec_1608;
  reg        [7:0]    regVec_1609;
  reg        [7:0]    regVec_1610;
  reg        [7:0]    regVec_1611;
  reg        [7:0]    regVec_1612;
  reg        [7:0]    regVec_1613;
  reg        [7:0]    regVec_1614;
  reg        [7:0]    regVec_1615;
  reg        [7:0]    regVec_1616;
  reg        [7:0]    regVec_1617;
  reg        [7:0]    regVec_1618;
  reg        [7:0]    regVec_1619;
  reg        [7:0]    regVec_1620;
  reg        [7:0]    regVec_1621;
  reg        [7:0]    regVec_1622;
  reg        [7:0]    regVec_1623;
  reg        [7:0]    regVec_1624;
  reg        [7:0]    regVec_1625;
  reg        [7:0]    regVec_1626;
  reg        [7:0]    regVec_1627;
  reg        [7:0]    regVec_1628;
  reg        [7:0]    regVec_1629;
  reg        [7:0]    regVec_1630;
  reg        [7:0]    regVec_1631;
  reg        [7:0]    regVec_1632;
  reg        [7:0]    regVec_1633;
  reg        [7:0]    regVec_1634;
  reg        [7:0]    regVec_1635;
  reg        [7:0]    regVec_1636;
  reg        [7:0]    regVec_1637;
  reg        [7:0]    regVec_1638;
  reg        [7:0]    regVec_1639;
  reg        [7:0]    regVec_1640;
  reg        [7:0]    regVec_1641;
  reg        [7:0]    regVec_1642;
  reg        [7:0]    regVec_1643;
  reg        [7:0]    regVec_1644;
  reg        [7:0]    regVec_1645;
  reg        [7:0]    regVec_1646;
  reg        [7:0]    regVec_1647;
  reg        [7:0]    regVec_1648;
  reg        [7:0]    regVec_1649;
  reg        [7:0]    regVec_1650;
  reg        [7:0]    regVec_1651;
  reg        [7:0]    regVec_1652;
  reg        [7:0]    regVec_1653;
  reg        [7:0]    regVec_1654;
  reg        [7:0]    regVec_1655;
  reg        [7:0]    regVec_1656;
  reg        [7:0]    regVec_1657;
  reg        [7:0]    regVec_1658;
  reg        [7:0]    regVec_1659;
  reg        [7:0]    regVec_1660;
  reg        [7:0]    regVec_1661;
  reg        [7:0]    regVec_1662;
  reg        [7:0]    regVec_1663;
  reg        [7:0]    regVec_1664;
  reg        [7:0]    regVec_1665;
  reg        [7:0]    regVec_1666;
  reg        [7:0]    regVec_1667;
  reg        [7:0]    regVec_1668;
  reg        [7:0]    regVec_1669;
  reg        [7:0]    regVec_1670;
  reg        [7:0]    regVec_1671;
  reg        [7:0]    regVec_1672;
  reg        [7:0]    regVec_1673;
  reg        [7:0]    regVec_1674;
  reg        [7:0]    regVec_1675;
  reg        [7:0]    regVec_1676;
  reg        [7:0]    regVec_1677;
  reg        [7:0]    regVec_1678;
  reg        [7:0]    regVec_1679;
  reg        [7:0]    regVec_1680;
  reg        [7:0]    regVec_1681;
  reg        [7:0]    regVec_1682;
  reg        [7:0]    regVec_1683;
  reg        [7:0]    regVec_1684;
  reg        [7:0]    regVec_1685;
  reg        [7:0]    regVec_1686;
  reg        [7:0]    regVec_1687;
  reg        [7:0]    regVec_1688;
  reg        [7:0]    regVec_1689;
  reg        [7:0]    regVec_1690;
  reg        [7:0]    regVec_1691;
  reg        [7:0]    regVec_1692;
  reg        [7:0]    regVec_1693;
  reg        [7:0]    regVec_1694;
  reg        [7:0]    regVec_1695;
  reg        [7:0]    regVec_1696;
  reg        [7:0]    regVec_1697;
  reg        [7:0]    regVec_1698;
  reg        [7:0]    regVec_1699;
  reg        [7:0]    regVec_1700;
  reg        [7:0]    regVec_1701;
  reg        [7:0]    regVec_1702;
  reg        [7:0]    regVec_1703;
  reg        [7:0]    regVec_1704;
  reg        [7:0]    regVec_1705;
  reg        [7:0]    regVec_1706;
  reg        [7:0]    regVec_1707;
  reg        [7:0]    regVec_1708;
  reg        [7:0]    regVec_1709;
  reg        [7:0]    regVec_1710;
  reg        [7:0]    regVec_1711;
  reg        [7:0]    regVec_1712;
  reg        [7:0]    regVec_1713;
  reg        [7:0]    regVec_1714;
  reg        [7:0]    regVec_1715;
  reg        [7:0]    regVec_1716;
  reg        [7:0]    regVec_1717;
  reg        [7:0]    regVec_1718;
  reg        [7:0]    regVec_1719;
  reg        [7:0]    regVec_1720;
  reg        [7:0]    regVec_1721;
  reg        [7:0]    regVec_1722;
  reg        [7:0]    regVec_1723;
  reg        [7:0]    regVec_1724;
  reg        [7:0]    regVec_1725;
  reg        [7:0]    regVec_1726;
  reg        [7:0]    regVec_1727;
  reg        [7:0]    regVec_1728;
  reg        [7:0]    regVec_1729;
  reg        [7:0]    regVec_1730;
  reg        [7:0]    regVec_1731;
  reg        [7:0]    regVec_1732;
  reg        [7:0]    regVec_1733;
  reg        [7:0]    regVec_1734;
  reg        [7:0]    regVec_1735;
  reg        [7:0]    regVec_1736;
  reg        [7:0]    regVec_1737;
  reg        [7:0]    regVec_1738;
  reg        [7:0]    regVec_1739;
  reg        [7:0]    regVec_1740;
  reg        [7:0]    regVec_1741;
  reg        [7:0]    regVec_1742;
  reg        [7:0]    regVec_1743;
  reg        [7:0]    regVec_1744;
  reg        [7:0]    regVec_1745;
  reg        [7:0]    regVec_1746;
  reg        [7:0]    regVec_1747;
  reg        [7:0]    regVec_1748;
  reg        [7:0]    regVec_1749;
  reg        [7:0]    regVec_1750;
  reg        [7:0]    regVec_1751;
  reg        [7:0]    regVec_1752;
  reg        [7:0]    regVec_1753;
  reg        [7:0]    regVec_1754;
  reg        [7:0]    regVec_1755;
  reg        [7:0]    regVec_1756;
  reg        [7:0]    regVec_1757;
  reg        [7:0]    regVec_1758;
  reg        [7:0]    regVec_1759;
  reg        [7:0]    regVec_1760;
  reg        [7:0]    regVec_1761;
  reg        [7:0]    regVec_1762;
  reg        [7:0]    regVec_1763;
  reg        [7:0]    regVec_1764;
  reg        [7:0]    regVec_1765;
  reg        [7:0]    regVec_1766;
  reg        [7:0]    regVec_1767;
  reg        [7:0]    regVec_1768;
  reg        [7:0]    regVec_1769;
  reg        [7:0]    regVec_1770;
  reg        [7:0]    regVec_1771;
  reg        [7:0]    regVec_1772;
  reg        [7:0]    regVec_1773;
  reg        [7:0]    regVec_1774;
  reg        [7:0]    regVec_1775;
  reg        [7:0]    regVec_1776;
  reg        [7:0]    regVec_1777;
  reg        [7:0]    regVec_1778;
  reg        [7:0]    regVec_1779;
  reg        [7:0]    regVec_1780;
  reg        [7:0]    regVec_1781;
  reg        [7:0]    regVec_1782;
  reg        [7:0]    regVec_1783;
  reg        [7:0]    regVec_1784;
  reg        [7:0]    regVec_1785;
  reg        [7:0]    regVec_1786;
  reg        [7:0]    regVec_1787;
  reg        [7:0]    regVec_1788;
  reg        [7:0]    regVec_1789;
  reg        [7:0]    regVec_1790;
  reg        [7:0]    regVec_1791;
  reg        [7:0]    regVec_1792;
  reg        [7:0]    regVec_1793;
  reg        [7:0]    regVec_1794;
  reg        [7:0]    regVec_1795;
  reg        [7:0]    regVec_1796;
  reg        [7:0]    regVec_1797;
  reg        [7:0]    regVec_1798;
  reg        [7:0]    regVec_1799;
  reg        [7:0]    regVec_1800;
  reg        [7:0]    regVec_1801;
  reg        [7:0]    regVec_1802;
  reg        [7:0]    regVec_1803;
  reg        [7:0]    regVec_1804;
  reg        [7:0]    regVec_1805;
  reg        [7:0]    regVec_1806;
  reg        [7:0]    regVec_1807;
  reg        [7:0]    regVec_1808;
  reg        [7:0]    regVec_1809;
  reg        [7:0]    regVec_1810;
  reg        [7:0]    regVec_1811;
  reg        [7:0]    regVec_1812;
  reg        [7:0]    regVec_1813;
  reg        [7:0]    regVec_1814;
  reg        [7:0]    regVec_1815;
  reg        [7:0]    regVec_1816;
  reg        [7:0]    regVec_1817;
  reg        [7:0]    regVec_1818;
  reg        [7:0]    regVec_1819;
  reg        [7:0]    regVec_1820;
  reg        [7:0]    regVec_1821;
  reg        [7:0]    regVec_1822;
  reg        [7:0]    regVec_1823;
  reg        [7:0]    regVec_1824;
  reg        [7:0]    regVec_1825;
  reg        [7:0]    regVec_1826;
  reg        [7:0]    regVec_1827;
  reg        [7:0]    regVec_1828;
  reg        [7:0]    regVec_1829;
  reg        [7:0]    regVec_1830;
  reg        [7:0]    regVec_1831;
  reg        [7:0]    regVec_1832;
  reg        [7:0]    regVec_1833;
  reg        [7:0]    regVec_1834;
  reg        [7:0]    regVec_1835;
  reg        [7:0]    regVec_1836;
  reg        [7:0]    regVec_1837;
  reg        [7:0]    regVec_1838;
  reg        [7:0]    regVec_1839;
  reg        [7:0]    regVec_1840;
  reg        [7:0]    regVec_1841;
  reg        [7:0]    regVec_1842;
  reg        [7:0]    regVec_1843;
  reg        [7:0]    regVec_1844;
  reg        [7:0]    regVec_1845;
  reg        [7:0]    regVec_1846;
  reg        [7:0]    regVec_1847;
  reg        [7:0]    regVec_1848;
  reg        [7:0]    regVec_1849;
  reg        [7:0]    regVec_1850;
  reg        [7:0]    regVec_1851;
  reg        [7:0]    regVec_1852;
  reg        [7:0]    regVec_1853;
  reg        [7:0]    regVec_1854;
  reg        [7:0]    regVec_1855;
  reg        [7:0]    regVec_1856;
  reg        [7:0]    regVec_1857;
  reg        [7:0]    regVec_1858;
  reg        [7:0]    regVec_1859;
  reg        [7:0]    regVec_1860;
  reg        [7:0]    regVec_1861;
  reg        [7:0]    regVec_1862;
  reg        [7:0]    regVec_1863;
  reg        [7:0]    regVec_1864;
  reg        [7:0]    regVec_1865;
  reg        [7:0]    regVec_1866;
  reg        [7:0]    regVec_1867;
  reg        [7:0]    regVec_1868;
  reg        [7:0]    regVec_1869;
  reg        [7:0]    regVec_1870;
  reg        [7:0]    regVec_1871;
  reg        [7:0]    regVec_1872;
  reg        [7:0]    regVec_1873;
  reg        [7:0]    regVec_1874;
  reg        [7:0]    regVec_1875;
  reg        [7:0]    regVec_1876;
  reg        [7:0]    regVec_1877;
  reg        [7:0]    regVec_1878;
  reg        [7:0]    regVec_1879;
  reg        [7:0]    regVec_1880;
  reg        [7:0]    regVec_1881;
  reg        [7:0]    regVec_1882;
  reg        [7:0]    regVec_1883;
  reg        [7:0]    regVec_1884;
  reg        [7:0]    regVec_1885;
  reg        [7:0]    regVec_1886;
  reg        [7:0]    regVec_1887;
  reg        [7:0]    regVec_1888;
  reg        [7:0]    regVec_1889;
  reg        [7:0]    regVec_1890;
  reg        [7:0]    regVec_1891;
  reg        [7:0]    regVec_1892;
  reg        [7:0]    regVec_1893;
  reg        [7:0]    regVec_1894;
  reg        [7:0]    regVec_1895;
  reg        [7:0]    regVec_1896;
  reg        [7:0]    regVec_1897;
  reg        [7:0]    regVec_1898;
  reg        [7:0]    regVec_1899;
  reg        [7:0]    regVec_1900;
  reg        [7:0]    regVec_1901;
  reg        [7:0]    regVec_1902;
  reg        [7:0]    regVec_1903;
  reg        [7:0]    regVec_1904;
  reg        [7:0]    regVec_1905;
  reg        [7:0]    regVec_1906;
  reg        [7:0]    regVec_1907;
  reg        [7:0]    regVec_1908;
  reg        [7:0]    regVec_1909;
  reg        [7:0]    regVec_1910;
  reg        [7:0]    regVec_1911;
  reg        [7:0]    regVec_1912;
  reg        [7:0]    regVec_1913;
  reg        [7:0]    regVec_1914;
  reg        [7:0]    regVec_1915;
  reg        [7:0]    regVec_1916;
  reg        [7:0]    regVec_1917;
  reg        [7:0]    regVec_1918;
  reg        [7:0]    regVec_1919;
  reg        [7:0]    regVec_1920;
  reg        [7:0]    regVec_1921;
  reg        [7:0]    regVec_1922;
  reg        [7:0]    regVec_1923;
  reg        [7:0]    regVec_1924;
  reg        [7:0]    regVec_1925;
  reg        [7:0]    regVec_1926;
  reg        [7:0]    regVec_1927;
  reg        [7:0]    regVec_1928;
  reg        [7:0]    regVec_1929;
  reg        [7:0]    regVec_1930;
  reg        [7:0]    regVec_1931;
  reg        [7:0]    regVec_1932;
  reg        [7:0]    regVec_1933;
  reg        [7:0]    regVec_1934;
  reg        [7:0]    regVec_1935;
  reg        [7:0]    regVec_1936;
  reg        [7:0]    regVec_1937;
  reg        [7:0]    regVec_1938;
  reg        [7:0]    regVec_1939;
  reg        [7:0]    regVec_1940;
  reg        [7:0]    regVec_1941;
  reg        [7:0]    regVec_1942;
  reg        [7:0]    regVec_1943;
  reg        [7:0]    regVec_1944;
  reg        [7:0]    regVec_1945;
  reg        [7:0]    regVec_1946;
  reg        [7:0]    regVec_1947;
  reg        [7:0]    regVec_1948;
  reg        [7:0]    regVec_1949;
  reg        [7:0]    regVec_1950;
  reg        [7:0]    regVec_1951;
  reg        [7:0]    regVec_1952;
  reg        [7:0]    regVec_1953;
  reg        [7:0]    regVec_1954;
  reg        [7:0]    regVec_1955;
  reg        [7:0]    regVec_1956;
  reg        [7:0]    regVec_1957;
  reg        [7:0]    regVec_1958;
  reg        [7:0]    regVec_1959;
  reg        [7:0]    regVec_1960;
  reg        [7:0]    regVec_1961;
  reg        [7:0]    regVec_1962;
  reg        [7:0]    regVec_1963;
  reg        [7:0]    regVec_1964;
  reg        [7:0]    regVec_1965;
  reg        [7:0]    regVec_1966;
  reg        [7:0]    regVec_1967;
  reg        [7:0]    regVec_1968;
  reg        [7:0]    regVec_1969;
  reg        [7:0]    regVec_1970;
  reg        [7:0]    regVec_1971;
  reg        [7:0]    regVec_1972;
  reg        [7:0]    regVec_1973;
  reg        [7:0]    regVec_1974;
  reg        [7:0]    regVec_1975;
  reg        [7:0]    regVec_1976;
  reg        [7:0]    regVec_1977;
  reg        [7:0]    regVec_1978;
  reg        [7:0]    regVec_1979;
  reg        [7:0]    regVec_1980;
  reg        [7:0]    regVec_1981;
  reg        [7:0]    regVec_1982;
  reg        [7:0]    regVec_1983;
  reg        [7:0]    regVec_1984;
  reg        [7:0]    regVec_1985;
  reg        [7:0]    regVec_1986;
  reg        [7:0]    regVec_1987;
  reg        [7:0]    regVec_1988;
  reg        [7:0]    regVec_1989;
  reg        [7:0]    regVec_1990;
  reg        [7:0]    regVec_1991;
  reg        [7:0]    regVec_1992;
  reg        [7:0]    regVec_1993;
  reg        [7:0]    regVec_1994;
  reg        [7:0]    regVec_1995;
  reg        [7:0]    regVec_1996;
  reg        [7:0]    regVec_1997;
  reg        [7:0]    regVec_1998;
  reg        [7:0]    regVec_1999;
  reg        [7:0]    regVec_2000;
  reg        [7:0]    regVec_2001;
  reg        [7:0]    regVec_2002;
  reg        [7:0]    regVec_2003;
  reg        [7:0]    regVec_2004;
  reg        [7:0]    regVec_2005;
  reg        [7:0]    regVec_2006;
  reg        [7:0]    regVec_2007;
  reg        [7:0]    regVec_2008;
  reg        [7:0]    regVec_2009;
  reg        [7:0]    regVec_2010;
  reg        [7:0]    regVec_2011;
  reg        [7:0]    regVec_2012;
  reg        [7:0]    regVec_2013;
  reg        [7:0]    regVec_2014;
  reg        [7:0]    regVec_2015;
  reg        [7:0]    regVec_2016;
  reg        [7:0]    regVec_2017;
  reg        [7:0]    regVec_2018;
  reg        [7:0]    regVec_2019;
  reg        [7:0]    regVec_2020;
  reg        [7:0]    regVec_2021;
  reg        [7:0]    regVec_2022;
  reg        [7:0]    regVec_2023;
  reg        [7:0]    regVec_2024;
  reg        [7:0]    regVec_2025;
  reg        [7:0]    regVec_2026;
  reg        [7:0]    regVec_2027;
  reg        [7:0]    regVec_2028;
  reg        [7:0]    regVec_2029;
  reg        [7:0]    regVec_2030;
  reg        [7:0]    regVec_2031;
  reg        [7:0]    regVec_2032;
  reg        [7:0]    regVec_2033;
  reg        [7:0]    regVec_2034;
  reg        [7:0]    regVec_2035;
  reg        [7:0]    regVec_2036;
  reg        [7:0]    regVec_2037;
  reg        [7:0]    regVec_2038;
  reg        [7:0]    regVec_2039;
  reg        [7:0]    regVec_2040;
  reg        [7:0]    regVec_2041;
  reg        [7:0]    regVec_2042;
  reg        [7:0]    regVec_2043;
  reg        [7:0]    regVec_2044;
  reg        [7:0]    regVec_2045;
  reg        [7:0]    regVec_2046;
  reg        [7:0]    regVec_2047;
  reg        [7:0]    regVec_2048;
  reg        [7:0]    regVec_2049;
  reg        [7:0]    regVec_2050;
  reg        [7:0]    regVec_2051;
  reg        [7:0]    regVec_2052;
  reg        [7:0]    regVec_2053;
  reg        [7:0]    regVec_2054;
  reg        [7:0]    regVec_2055;
  reg        [7:0]    regVec_2056;
  reg        [7:0]    regVec_2057;
  reg        [7:0]    regVec_2058;
  reg        [7:0]    regVec_2059;
  reg        [7:0]    regVec_2060;
  reg        [7:0]    regVec_2061;
  reg        [7:0]    regVec_2062;
  reg        [7:0]    regVec_2063;
  reg        [7:0]    regVec_2064;
  reg        [7:0]    regVec_2065;
  reg        [7:0]    regVec_2066;
  reg        [7:0]    regVec_2067;
  reg        [7:0]    regVec_2068;
  reg        [7:0]    regVec_2069;
  reg        [7:0]    regVec_2070;
  reg        [7:0]    regVec_2071;
  reg        [7:0]    regVec_2072;
  reg        [7:0]    regVec_2073;
  reg        [7:0]    regVec_2074;
  reg        [7:0]    regVec_2075;
  reg        [7:0]    regVec_2076;
  reg        [7:0]    regVec_2077;
  reg        [7:0]    regVec_2078;
  reg        [7:0]    regVec_2079;
  reg        [7:0]    regVec_2080;
  reg        [7:0]    regVec_2081;
  reg        [7:0]    regVec_2082;
  reg        [7:0]    regVec_2083;
  reg        [7:0]    regVec_2084;
  reg        [7:0]    regVec_2085;
  reg        [7:0]    regVec_2086;
  reg        [7:0]    regVec_2087;
  reg        [7:0]    regVec_2088;
  reg        [7:0]    regVec_2089;
  reg        [7:0]    regVec_2090;
  reg        [7:0]    regVec_2091;
  reg        [7:0]    regVec_2092;
  reg        [7:0]    regVec_2093;
  reg        [7:0]    regVec_2094;
  reg        [7:0]    regVec_2095;
  reg        [7:0]    regVec_2096;
  reg        [7:0]    regVec_2097;
  reg        [7:0]    regVec_2098;
  reg        [7:0]    regVec_2099;
  reg        [7:0]    regVec_2100;
  reg        [7:0]    regVec_2101;
  reg        [7:0]    regVec_2102;
  reg        [7:0]    regVec_2103;
  reg        [7:0]    regVec_2104;
  reg        [7:0]    regVec_2105;
  reg        [7:0]    regVec_2106;
  reg        [7:0]    regVec_2107;
  reg        [7:0]    regVec_2108;
  reg        [7:0]    regVec_2109;
  reg        [7:0]    regVec_2110;
  reg        [7:0]    regVec_2111;
  reg        [7:0]    regVec_2112;
  reg        [7:0]    regVec_2113;
  reg        [7:0]    regVec_2114;
  reg        [7:0]    regVec_2115;
  reg        [7:0]    regVec_2116;
  reg        [7:0]    regVec_2117;
  reg        [7:0]    regVec_2118;
  reg        [7:0]    regVec_2119;
  reg        [7:0]    regVec_2120;
  reg        [7:0]    regVec_2121;
  reg        [7:0]    regVec_2122;
  reg        [7:0]    regVec_2123;
  reg        [7:0]    regVec_2124;
  reg        [7:0]    regVec_2125;
  reg        [7:0]    regVec_2126;
  reg        [7:0]    regVec_2127;
  reg        [7:0]    regVec_2128;
  reg        [7:0]    regVec_2129;
  reg        [7:0]    regVec_2130;
  reg        [7:0]    regVec_2131;
  reg        [7:0]    regVec_2132;
  reg        [7:0]    regVec_2133;
  reg        [7:0]    regVec_2134;
  reg        [7:0]    regVec_2135;
  reg        [7:0]    regVec_2136;
  reg        [7:0]    regVec_2137;
  reg        [7:0]    regVec_2138;
  reg        [7:0]    regVec_2139;
  reg        [7:0]    regVec_2140;
  reg        [7:0]    regVec_2141;
  reg        [7:0]    regVec_2142;
  reg        [7:0]    regVec_2143;
  reg        [7:0]    regVec_2144;
  reg        [7:0]    regVec_2145;
  reg        [7:0]    regVec_2146;
  reg        [7:0]    regVec_2147;
  reg        [7:0]    regVec_2148;
  reg        [7:0]    regVec_2149;
  reg        [7:0]    regVec_2150;
  reg        [7:0]    regVec_2151;
  reg        [7:0]    regVec_2152;
  reg        [7:0]    regVec_2153;
  reg        [7:0]    regVec_2154;
  reg        [7:0]    regVec_2155;
  reg        [7:0]    regVec_2156;
  reg        [7:0]    regVec_2157;
  reg        [7:0]    regVec_2158;
  reg        [7:0]    regVec_2159;
  reg        [7:0]    regVec_2160;
  reg        [7:0]    regVec_2161;
  reg        [7:0]    regVec_2162;
  reg        [7:0]    regVec_2163;
  reg        [7:0]    regVec_2164;
  reg        [7:0]    regVec_2165;
  reg        [7:0]    regVec_2166;
  reg        [7:0]    regVec_2167;
  reg        [7:0]    regVec_2168;
  reg        [7:0]    regVec_2169;
  reg        [7:0]    regVec_2170;
  reg        [7:0]    regVec_2171;
  reg        [7:0]    regVec_2172;
  reg        [7:0]    regVec_2173;
  reg        [7:0]    regVec_2174;
  reg        [7:0]    regVec_2175;
  reg        [7:0]    regVec_2176;
  reg        [7:0]    regVec_2177;
  reg        [7:0]    regVec_2178;
  reg        [7:0]    regVec_2179;
  reg        [7:0]    regVec_2180;
  reg        [7:0]    regVec_2181;
  reg        [7:0]    regVec_2182;
  reg        [7:0]    regVec_2183;
  reg        [7:0]    regVec_2184;
  reg        [7:0]    regVec_2185;
  reg        [7:0]    regVec_2186;
  reg        [7:0]    regVec_2187;
  reg        [7:0]    regVec_2188;
  reg        [7:0]    regVec_2189;
  reg        [7:0]    regVec_2190;
  reg        [7:0]    regVec_2191;
  reg        [7:0]    regVec_2192;
  reg        [7:0]    regVec_2193;
  reg        [7:0]    regVec_2194;
  reg        [7:0]    regVec_2195;
  reg        [7:0]    regVec_2196;
  reg        [7:0]    regVec_2197;
  reg        [7:0]    regVec_2198;
  reg        [7:0]    regVec_2199;
  reg        [7:0]    regVec_2200;
  reg        [7:0]    regVec_2201;
  reg        [7:0]    regVec_2202;
  reg        [7:0]    regVec_2203;
  reg        [7:0]    regVec_2204;
  reg        [7:0]    regVec_2205;
  reg        [7:0]    regVec_2206;
  reg        [7:0]    regVec_2207;
  reg        [7:0]    regVec_2208;
  reg        [7:0]    regVec_2209;
  reg        [7:0]    regVec_2210;
  reg        [7:0]    regVec_2211;
  reg        [7:0]    regVec_2212;
  reg        [7:0]    regVec_2213;
  reg        [7:0]    regVec_2214;
  reg        [7:0]    regVec_2215;
  reg        [7:0]    regVec_2216;
  reg        [7:0]    regVec_2217;
  reg        [7:0]    regVec_2218;
  reg        [7:0]    regVec_2219;
  reg        [7:0]    regVec_2220;
  reg        [7:0]    regVec_2221;
  reg        [7:0]    regVec_2222;
  reg        [7:0]    regVec_2223;
  reg        [7:0]    regVec_2224;
  reg        [7:0]    regVec_2225;
  reg        [7:0]    regVec_2226;
  reg        [7:0]    regVec_2227;
  reg        [7:0]    regVec_2228;
  reg        [7:0]    regVec_2229;
  reg        [7:0]    regVec_2230;
  reg        [7:0]    regVec_2231;
  reg        [7:0]    regVec_2232;
  reg        [7:0]    regVec_2233;
  reg        [7:0]    regVec_2234;
  reg        [7:0]    regVec_2235;
  reg        [7:0]    regVec_2236;
  reg        [7:0]    regVec_2237;
  reg        [7:0]    regVec_2238;
  reg        [7:0]    regVec_2239;
  reg        [7:0]    regVec_2240;
  reg        [7:0]    regVec_2241;
  reg        [7:0]    regVec_2242;
  reg        [7:0]    regVec_2243;
  reg        [7:0]    regVec_2244;
  reg        [7:0]    regVec_2245;
  reg        [7:0]    regVec_2246;
  reg        [7:0]    regVec_2247;
  reg        [7:0]    regVec_2248;
  reg        [7:0]    regVec_2249;
  reg        [7:0]    regVec_2250;
  reg        [7:0]    regVec_2251;
  reg        [7:0]    regVec_2252;
  reg        [7:0]    regVec_2253;
  reg        [7:0]    regVec_2254;
  reg        [7:0]    regVec_2255;
  reg        [7:0]    regVec_2256;
  reg        [7:0]    regVec_2257;
  reg        [7:0]    regVec_2258;
  reg        [7:0]    regVec_2259;
  reg        [7:0]    regVec_2260;
  reg        [7:0]    regVec_2261;
  reg        [7:0]    regVec_2262;
  reg        [7:0]    regVec_2263;
  reg        [7:0]    regVec_2264;
  reg        [7:0]    regVec_2265;
  reg        [7:0]    regVec_2266;
  reg        [7:0]    regVec_2267;
  reg        [7:0]    regVec_2268;
  reg        [7:0]    regVec_2269;
  reg        [7:0]    regVec_2270;
  reg        [7:0]    regVec_2271;
  reg        [7:0]    regVec_2272;
  reg        [7:0]    regVec_2273;
  reg        [7:0]    regVec_2274;
  reg        [7:0]    regVec_2275;
  reg        [7:0]    regVec_2276;
  reg        [7:0]    regVec_2277;
  reg        [7:0]    regVec_2278;
  reg        [7:0]    regVec_2279;
  reg        [7:0]    regVec_2280;
  reg        [7:0]    regVec_2281;
  reg        [7:0]    regVec_2282;
  reg        [7:0]    regVec_2283;
  reg        [7:0]    regVec_2284;
  reg        [7:0]    regVec_2285;
  reg        [7:0]    regVec_2286;
  reg        [7:0]    regVec_2287;
  reg        [7:0]    regVec_2288;
  reg        [7:0]    regVec_2289;
  reg        [7:0]    regVec_2290;
  reg        [7:0]    regVec_2291;
  reg        [7:0]    regVec_2292;
  reg        [7:0]    regVec_2293;
  reg        [7:0]    regVec_2294;
  reg        [7:0]    regVec_2295;
  reg        [7:0]    regVec_2296;
  reg        [7:0]    regVec_2297;
  reg        [7:0]    regVec_2298;
  reg        [7:0]    regVec_2299;
  reg        [7:0]    regVec_2300;
  reg        [7:0]    regVec_2301;
  reg        [7:0]    regVec_2302;
  reg        [7:0]    regVec_2303;
  reg        [7:0]    regVec_2304;
  reg        [7:0]    regVec_2305;
  reg        [7:0]    regVec_2306;
  reg        [7:0]    regVec_2307;
  reg        [7:0]    regVec_2308;
  reg        [7:0]    regVec_2309;
  reg        [7:0]    regVec_2310;
  reg        [7:0]    regVec_2311;
  reg        [7:0]    regVec_2312;
  reg        [7:0]    regVec_2313;
  reg        [7:0]    regVec_2314;
  reg        [7:0]    regVec_2315;
  reg        [7:0]    regVec_2316;
  reg        [7:0]    regVec_2317;
  reg        [7:0]    regVec_2318;
  reg        [7:0]    regVec_2319;
  reg        [7:0]    regVec_2320;
  reg        [7:0]    regVec_2321;
  reg        [7:0]    regVec_2322;
  reg        [7:0]    regVec_2323;
  reg        [7:0]    regVec_2324;
  reg        [7:0]    regVec_2325;
  reg        [7:0]    regVec_2326;
  reg        [7:0]    regVec_2327;
  reg        [7:0]    regVec_2328;
  reg        [7:0]    regVec_2329;
  reg        [7:0]    regVec_2330;
  reg        [7:0]    regVec_2331;
  reg        [7:0]    regVec_2332;
  reg        [7:0]    regVec_2333;
  reg        [7:0]    regVec_2334;
  reg        [7:0]    regVec_2335;
  reg        [7:0]    regVec_2336;
  reg        [7:0]    regVec_2337;
  reg        [7:0]    regVec_2338;
  reg        [7:0]    regVec_2339;
  reg        [7:0]    regVec_2340;
  reg        [7:0]    regVec_2341;
  reg        [7:0]    regVec_2342;
  reg        [7:0]    regVec_2343;
  reg        [7:0]    regVec_2344;
  reg        [7:0]    regVec_2345;
  reg        [7:0]    regVec_2346;
  reg        [7:0]    regVec_2347;
  reg        [7:0]    regVec_2348;
  reg        [7:0]    regVec_2349;
  reg        [7:0]    regVec_2350;
  reg        [7:0]    regVec_2351;
  reg        [7:0]    regVec_2352;
  reg        [7:0]    regVec_2353;
  reg        [7:0]    regVec_2354;
  reg        [7:0]    regVec_2355;
  reg        [7:0]    regVec_2356;
  reg        [7:0]    regVec_2357;
  reg        [7:0]    regVec_2358;
  reg        [7:0]    regVec_2359;
  reg        [7:0]    regVec_2360;
  reg        [7:0]    regVec_2361;
  reg        [7:0]    regVec_2362;
  reg        [7:0]    regVec_2363;
  reg        [7:0]    regVec_2364;
  reg        [7:0]    regVec_2365;
  reg        [7:0]    regVec_2366;
  reg        [7:0]    regVec_2367;
  reg        [7:0]    regVec_2368;
  reg        [7:0]    regVec_2369;
  reg        [7:0]    regVec_2370;
  reg        [7:0]    regVec_2371;
  reg        [7:0]    regVec_2372;
  reg        [7:0]    regVec_2373;
  reg        [7:0]    regVec_2374;
  reg        [7:0]    regVec_2375;
  reg        [7:0]    regVec_2376;
  reg        [7:0]    regVec_2377;
  reg        [7:0]    regVec_2378;
  reg        [7:0]    regVec_2379;
  reg        [7:0]    regVec_2380;
  reg        [7:0]    regVec_2381;
  reg        [7:0]    regVec_2382;
  reg        [7:0]    regVec_2383;
  reg        [7:0]    regVec_2384;
  reg        [7:0]    regVec_2385;
  reg        [7:0]    regVec_2386;
  reg        [7:0]    regVec_2387;
  reg        [7:0]    regVec_2388;
  reg        [7:0]    regVec_2389;
  reg        [7:0]    regVec_2390;
  reg        [7:0]    regVec_2391;
  reg        [7:0]    regVec_2392;
  reg        [7:0]    regVec_2393;
  reg        [7:0]    regVec_2394;
  reg        [7:0]    regVec_2395;
  reg        [7:0]    regVec_2396;
  reg        [7:0]    regVec_2397;
  reg        [7:0]    regVec_2398;
  reg        [7:0]    regVec_2399;
  reg        [7:0]    regVec_2400;
  reg        [7:0]    regVec_2401;
  reg        [7:0]    regVec_2402;
  reg        [7:0]    regVec_2403;
  reg        [7:0]    regVec_2404;
  reg        [7:0]    regVec_2405;
  reg        [7:0]    regVec_2406;
  reg        [7:0]    regVec_2407;
  reg        [7:0]    regVec_2408;
  reg        [7:0]    regVec_2409;
  reg        [7:0]    regVec_2410;
  reg        [7:0]    regVec_2411;
  reg        [7:0]    regVec_2412;
  reg        [7:0]    regVec_2413;
  reg        [7:0]    regVec_2414;
  reg        [7:0]    regVec_2415;
  reg        [7:0]    regVec_2416;
  reg        [7:0]    regVec_2417;
  reg        [7:0]    regVec_2418;
  reg        [7:0]    regVec_2419;
  reg        [7:0]    regVec_2420;
  reg        [7:0]    regVec_2421;
  reg        [7:0]    regVec_2422;
  reg        [7:0]    regVec_2423;
  reg        [7:0]    regVec_2424;
  reg        [7:0]    regVec_2425;
  reg        [7:0]    regVec_2426;
  reg        [7:0]    regVec_2427;
  reg        [7:0]    regVec_2428;
  reg        [7:0]    regVec_2429;
  reg        [7:0]    regVec_2430;
  reg        [7:0]    regVec_2431;
  reg        [7:0]    regVec_2432;
  reg        [7:0]    regVec_2433;
  reg        [7:0]    regVec_2434;
  reg        [7:0]    regVec_2435;
  reg        [7:0]    regVec_2436;
  reg        [7:0]    regVec_2437;
  reg        [7:0]    regVec_2438;
  reg        [7:0]    regVec_2439;
  reg        [7:0]    regVec_2440;
  reg        [7:0]    regVec_2441;
  reg        [7:0]    regVec_2442;
  reg        [7:0]    regVec_2443;
  reg        [7:0]    regVec_2444;
  reg        [7:0]    regVec_2445;
  reg        [7:0]    regVec_2446;
  reg        [7:0]    regVec_2447;
  reg        [7:0]    regVec_2448;
  reg        [7:0]    regVec_2449;
  reg        [7:0]    regVec_2450;
  reg        [7:0]    regVec_2451;
  reg        [7:0]    regVec_2452;
  reg        [7:0]    regVec_2453;
  reg        [7:0]    regVec_2454;
  reg        [7:0]    regVec_2455;
  reg        [7:0]    regVec_2456;
  reg        [7:0]    regVec_2457;
  reg        [7:0]    regVec_2458;
  reg        [7:0]    regVec_2459;
  reg        [7:0]    regVec_2460;
  reg        [7:0]    regVec_2461;
  reg        [7:0]    regVec_2462;
  reg        [7:0]    regVec_2463;
  reg        [7:0]    regVec_2464;
  reg        [7:0]    regVec_2465;
  reg        [7:0]    regVec_2466;
  reg        [7:0]    regVec_2467;
  reg        [7:0]    regVec_2468;
  reg        [7:0]    regVec_2469;
  reg        [7:0]    regVec_2470;
  reg        [7:0]    regVec_2471;
  reg        [7:0]    regVec_2472;
  reg        [7:0]    regVec_2473;
  reg        [7:0]    regVec_2474;
  reg        [7:0]    regVec_2475;
  reg        [7:0]    regVec_2476;
  reg        [7:0]    regVec_2477;
  reg        [7:0]    regVec_2478;
  reg        [7:0]    regVec_2479;
  reg        [7:0]    regVec_2480;
  reg        [7:0]    regVec_2481;
  reg        [7:0]    regVec_2482;
  reg        [7:0]    regVec_2483;
  reg        [7:0]    regVec_2484;
  reg        [7:0]    regVec_2485;
  reg        [7:0]    regVec_2486;
  reg        [7:0]    regVec_2487;
  reg        [7:0]    regVec_2488;
  reg        [7:0]    regVec_2489;
  reg        [7:0]    regVec_2490;
  reg        [7:0]    regVec_2491;
  reg        [7:0]    regVec_2492;
  reg        [7:0]    regVec_2493;
  reg        [7:0]    regVec_2494;
  reg        [7:0]    regVec_2495;
  reg        [7:0]    regVec_2496;
  reg        [7:0]    regVec_2497;
  reg        [7:0]    regVec_2498;
  reg        [7:0]    regVec_2499;
  reg        [7:0]    regVec_2500;
  reg        [7:0]    regVec_2501;
  reg        [7:0]    regVec_2502;
  reg        [7:0]    regVec_2503;
  reg        [7:0]    regVec_2504;
  reg        [7:0]    regVec_2505;
  reg        [7:0]    regVec_2506;
  reg        [7:0]    regVec_2507;
  reg        [7:0]    regVec_2508;
  reg        [7:0]    regVec_2509;
  reg        [7:0]    regVec_2510;
  reg        [7:0]    regVec_2511;
  reg        [7:0]    regVec_2512;
  reg        [7:0]    regVec_2513;
  reg        [7:0]    regVec_2514;
  reg        [7:0]    regVec_2515;
  reg        [7:0]    regVec_2516;
  reg        [7:0]    regVec_2517;
  reg        [7:0]    regVec_2518;
  reg        [7:0]    regVec_2519;
  reg        [7:0]    regVec_2520;
  reg        [7:0]    regVec_2521;
  reg        [7:0]    regVec_2522;
  reg        [7:0]    regVec_2523;
  reg        [7:0]    regVec_2524;
  reg        [7:0]    regVec_2525;
  reg        [7:0]    regVec_2526;
  reg        [7:0]    regVec_2527;
  reg        [7:0]    regVec_2528;
  reg        [7:0]    regVec_2529;
  reg        [7:0]    regVec_2530;
  reg        [7:0]    regVec_2531;
  reg        [7:0]    regVec_2532;
  reg        [7:0]    regVec_2533;
  reg        [7:0]    regVec_2534;
  reg        [7:0]    regVec_2535;
  reg        [7:0]    regVec_2536;
  reg        [7:0]    regVec_2537;
  reg        [7:0]    regVec_2538;
  reg        [7:0]    regVec_2539;
  reg        [7:0]    regVec_2540;
  reg        [7:0]    regVec_2541;
  reg        [7:0]    regVec_2542;
  reg        [7:0]    regVec_2543;
  reg        [7:0]    regVec_2544;
  reg        [7:0]    regVec_2545;
  reg        [7:0]    regVec_2546;
  reg        [7:0]    regVec_2547;
  reg        [7:0]    regVec_2548;
  reg        [7:0]    regVec_2549;
  reg        [7:0]    regVec_2550;
  reg        [7:0]    regVec_2551;
  reg        [7:0]    regVec_2552;
  reg        [7:0]    regVec_2553;
  reg        [7:0]    regVec_2554;
  reg        [7:0]    regVec_2555;
  reg        [7:0]    regVec_2556;
  reg        [7:0]    regVec_2557;
  reg        [7:0]    regVec_2558;
  reg        [7:0]    regVec_2559;
  reg        [7:0]    regVec_2560;
  reg        [7:0]    regVec_2561;
  reg        [7:0]    regVec_2562;
  reg        [7:0]    regVec_2563;
  reg        [7:0]    regVec_2564;
  reg        [7:0]    regVec_2565;
  reg        [7:0]    regVec_2566;
  reg        [7:0]    regVec_2567;
  reg        [7:0]    regVec_2568;
  reg        [7:0]    regVec_2569;
  reg        [7:0]    regVec_2570;
  reg        [7:0]    regVec_2571;
  reg        [7:0]    regVec_2572;
  reg        [7:0]    regVec_2573;
  reg        [7:0]    regVec_2574;
  reg        [7:0]    regVec_2575;
  reg        [7:0]    regVec_2576;
  reg        [7:0]    regVec_2577;
  reg        [7:0]    regVec_2578;
  reg        [7:0]    regVec_2579;
  reg        [7:0]    regVec_2580;
  reg        [7:0]    regVec_2581;
  reg        [7:0]    regVec_2582;
  reg        [7:0]    regVec_2583;
  reg        [7:0]    regVec_2584;
  reg        [7:0]    regVec_2585;
  reg        [7:0]    regVec_2586;
  reg        [7:0]    regVec_2587;
  reg        [7:0]    regVec_2588;
  reg        [7:0]    regVec_2589;
  reg        [7:0]    regVec_2590;
  reg        [7:0]    regVec_2591;
  reg        [7:0]    regVec_2592;
  reg        [7:0]    regVec_2593;
  reg        [7:0]    regVec_2594;
  reg        [7:0]    regVec_2595;
  reg        [7:0]    regVec_2596;
  reg        [7:0]    regVec_2597;
  reg        [7:0]    regVec_2598;
  reg        [7:0]    regVec_2599;
  reg        [7:0]    regVec_2600;
  reg        [7:0]    regVec_2601;
  reg        [7:0]    regVec_2602;
  reg        [7:0]    regVec_2603;
  reg        [7:0]    regVec_2604;
  reg        [7:0]    regVec_2605;
  reg        [7:0]    regVec_2606;
  reg        [7:0]    regVec_2607;
  reg        [7:0]    regVec_2608;
  reg        [7:0]    regVec_2609;
  reg        [7:0]    regVec_2610;
  reg        [7:0]    regVec_2611;
  reg        [7:0]    regVec_2612;
  reg        [7:0]    regVec_2613;
  reg        [7:0]    regVec_2614;
  reg        [7:0]    regVec_2615;
  reg        [7:0]    regVec_2616;
  reg        [7:0]    regVec_2617;
  reg        [7:0]    regVec_2618;
  reg        [7:0]    regVec_2619;
  reg        [7:0]    regVec_2620;
  reg        [7:0]    regVec_2621;
  reg        [7:0]    regVec_2622;
  reg        [7:0]    regVec_2623;
  reg        [7:0]    regVec_2624;
  reg        [7:0]    regVec_2625;
  reg        [7:0]    regVec_2626;
  reg        [7:0]    regVec_2627;
  reg        [7:0]    regVec_2628;
  reg        [7:0]    regVec_2629;
  reg        [7:0]    regVec_2630;
  reg        [7:0]    regVec_2631;
  reg        [7:0]    regVec_2632;
  reg        [7:0]    regVec_2633;
  reg        [7:0]    regVec_2634;
  reg        [7:0]    regVec_2635;
  reg        [7:0]    regVec_2636;
  reg        [7:0]    regVec_2637;
  reg        [7:0]    regVec_2638;
  reg        [7:0]    regVec_2639;
  reg        [7:0]    regVec_2640;
  reg        [7:0]    regVec_2641;
  reg        [7:0]    regVec_2642;
  reg        [7:0]    regVec_2643;
  reg        [7:0]    regVec_2644;
  reg        [7:0]    regVec_2645;
  reg        [7:0]    regVec_2646;
  reg        [7:0]    regVec_2647;
  reg        [7:0]    regVec_2648;
  reg        [7:0]    regVec_2649;
  reg        [7:0]    regVec_2650;
  reg        [7:0]    regVec_2651;
  reg        [7:0]    regVec_2652;
  reg        [7:0]    regVec_2653;
  reg        [7:0]    regVec_2654;
  reg        [7:0]    regVec_2655;
  reg        [7:0]    regVec_2656;
  reg        [7:0]    regVec_2657;
  reg        [7:0]    regVec_2658;
  reg        [7:0]    regVec_2659;
  reg        [7:0]    regVec_2660;
  reg        [7:0]    regVec_2661;
  reg        [7:0]    regVec_2662;
  reg        [7:0]    regVec_2663;
  reg        [7:0]    regVec_2664;
  reg        [7:0]    regVec_2665;
  reg        [7:0]    regVec_2666;
  reg        [7:0]    regVec_2667;
  reg        [7:0]    regVec_2668;
  reg        [7:0]    regVec_2669;
  reg        [7:0]    regVec_2670;
  reg        [7:0]    regVec_2671;
  reg        [7:0]    regVec_2672;
  reg        [7:0]    regVec_2673;
  reg        [7:0]    regVec_2674;
  reg        [7:0]    regVec_2675;
  reg        [7:0]    regVec_2676;
  reg        [7:0]    regVec_2677;
  reg        [7:0]    regVec_2678;
  reg        [7:0]    regVec_2679;
  reg        [7:0]    regVec_2680;
  reg        [7:0]    regVec_2681;
  reg        [7:0]    regVec_2682;
  reg        [7:0]    regVec_2683;
  reg        [7:0]    regVec_2684;
  reg        [7:0]    regVec_2685;
  reg        [7:0]    regVec_2686;
  reg        [7:0]    regVec_2687;
  reg        [7:0]    regVec_2688;
  reg        [7:0]    regVec_2689;
  reg        [7:0]    regVec_2690;
  reg        [7:0]    regVec_2691;
  reg        [7:0]    regVec_2692;
  reg        [7:0]    regVec_2693;
  reg        [7:0]    regVec_2694;
  reg        [7:0]    regVec_2695;
  reg        [7:0]    regVec_2696;
  reg        [7:0]    regVec_2697;
  reg        [7:0]    regVec_2698;
  reg        [7:0]    regVec_2699;
  reg        [7:0]    regVec_2700;
  reg        [7:0]    regVec_2701;
  reg        [7:0]    regVec_2702;
  reg        [7:0]    regVec_2703;
  reg        [7:0]    regVec_2704;
  reg        [7:0]    regVec_2705;
  reg        [7:0]    regVec_2706;
  reg        [7:0]    regVec_2707;
  reg        [7:0]    regVec_2708;
  reg        [7:0]    regVec_2709;
  reg        [7:0]    regVec_2710;
  reg        [7:0]    regVec_2711;
  reg        [7:0]    regVec_2712;
  reg        [7:0]    regVec_2713;
  reg        [7:0]    regVec_2714;
  reg        [7:0]    regVec_2715;
  reg        [7:0]    regVec_2716;
  reg        [7:0]    regVec_2717;
  reg        [7:0]    regVec_2718;
  reg        [7:0]    regVec_2719;
  reg        [7:0]    regVec_2720;
  reg        [7:0]    regVec_2721;
  reg        [7:0]    regVec_2722;
  reg        [7:0]    regVec_2723;
  reg        [7:0]    regVec_2724;
  reg        [7:0]    regVec_2725;
  reg        [7:0]    regVec_2726;
  reg        [7:0]    regVec_2727;
  reg        [7:0]    regVec_2728;
  reg        [7:0]    regVec_2729;
  reg        [7:0]    regVec_2730;
  reg        [7:0]    regVec_2731;
  reg        [7:0]    regVec_2732;
  reg        [7:0]    regVec_2733;
  reg        [7:0]    regVec_2734;
  reg        [7:0]    regVec_2735;
  reg        [7:0]    regVec_2736;
  reg        [7:0]    regVec_2737;
  reg        [7:0]    regVec_2738;
  reg        [7:0]    regVec_2739;
  reg        [7:0]    regVec_2740;
  reg        [7:0]    regVec_2741;
  reg        [7:0]    regVec_2742;
  reg        [7:0]    regVec_2743;
  reg        [7:0]    regVec_2744;
  reg        [7:0]    regVec_2745;
  reg        [7:0]    regVec_2746;
  reg        [7:0]    regVec_2747;
  reg        [7:0]    regVec_2748;
  reg        [7:0]    regVec_2749;
  reg        [7:0]    regVec_2750;
  reg        [7:0]    regVec_2751;
  reg        [7:0]    regVec_2752;
  reg        [7:0]    regVec_2753;
  reg        [7:0]    regVec_2754;
  reg        [7:0]    regVec_2755;
  reg        [7:0]    regVec_2756;
  reg        [7:0]    regVec_2757;
  reg        [7:0]    regVec_2758;
  reg        [7:0]    regVec_2759;
  reg        [7:0]    regVec_2760;
  reg        [7:0]    regVec_2761;
  reg        [7:0]    regVec_2762;
  reg        [7:0]    regVec_2763;
  reg        [7:0]    regVec_2764;
  reg        [7:0]    regVec_2765;
  reg        [7:0]    regVec_2766;
  reg        [7:0]    regVec_2767;
  reg        [7:0]    regVec_2768;
  reg        [7:0]    regVec_2769;
  reg        [7:0]    regVec_2770;
  reg        [7:0]    regVec_2771;
  reg        [7:0]    regVec_2772;
  reg        [7:0]    regVec_2773;
  reg        [7:0]    regVec_2774;
  reg        [7:0]    regVec_2775;
  reg        [7:0]    regVec_2776;
  reg        [7:0]    regVec_2777;
  reg        [7:0]    regVec_2778;
  reg        [7:0]    regVec_2779;
  reg        [7:0]    regVec_2780;
  reg        [7:0]    regVec_2781;
  reg        [7:0]    regVec_2782;
  reg        [7:0]    regVec_2783;
  reg        [7:0]    regVec_2784;
  reg        [7:0]    regVec_2785;
  reg        [7:0]    regVec_2786;
  reg        [7:0]    regVec_2787;
  reg        [7:0]    regVec_2788;
  reg        [7:0]    regVec_2789;
  reg        [7:0]    regVec_2790;
  reg        [7:0]    regVec_2791;
  reg        [7:0]    regVec_2792;
  reg        [7:0]    regVec_2793;
  reg        [7:0]    regVec_2794;
  reg        [7:0]    regVec_2795;
  reg        [7:0]    regVec_2796;
  reg        [7:0]    regVec_2797;
  reg        [7:0]    regVec_2798;
  reg        [7:0]    regVec_2799;
  reg        [7:0]    regVec_2800;
  reg        [7:0]    regVec_2801;
  reg        [7:0]    regVec_2802;
  reg        [7:0]    regVec_2803;
  reg        [7:0]    regVec_2804;
  reg        [7:0]    regVec_2805;
  reg        [7:0]    regVec_2806;
  reg        [7:0]    regVec_2807;
  reg        [7:0]    regVec_2808;
  reg        [7:0]    regVec_2809;
  reg        [7:0]    regVec_2810;
  reg        [7:0]    regVec_2811;
  reg        [7:0]    regVec_2812;
  reg        [7:0]    regVec_2813;
  reg        [7:0]    regVec_2814;
  reg        [7:0]    regVec_2815;
  reg        [7:0]    regVec_2816;
  reg        [7:0]    regVec_2817;
  reg        [7:0]    regVec_2818;
  reg        [7:0]    regVec_2819;
  reg        [7:0]    regVec_2820;
  reg        [7:0]    regVec_2821;
  reg        [7:0]    regVec_2822;
  reg        [7:0]    regVec_2823;
  reg        [7:0]    regVec_2824;
  reg        [7:0]    regVec_2825;
  reg        [7:0]    regVec_2826;
  reg        [7:0]    regVec_2827;
  reg        [7:0]    regVec_2828;
  reg        [7:0]    regVec_2829;
  reg        [7:0]    regVec_2830;
  reg        [7:0]    regVec_2831;
  reg        [7:0]    regVec_2832;
  reg        [7:0]    regVec_2833;
  reg        [7:0]    regVec_2834;
  reg        [7:0]    regVec_2835;
  reg        [7:0]    regVec_2836;
  reg        [7:0]    regVec_2837;
  reg        [7:0]    regVec_2838;
  reg        [7:0]    regVec_2839;
  reg        [7:0]    regVec_2840;
  reg        [7:0]    regVec_2841;
  reg        [7:0]    regVec_2842;
  reg        [7:0]    regVec_2843;
  reg        [7:0]    regVec_2844;
  reg        [7:0]    regVec_2845;
  reg        [7:0]    regVec_2846;
  reg        [7:0]    regVec_2847;
  reg        [7:0]    regVec_2848;
  reg        [7:0]    regVec_2849;
  reg        [7:0]    regVec_2850;
  reg        [7:0]    regVec_2851;
  reg        [7:0]    regVec_2852;
  reg        [7:0]    regVec_2853;
  reg        [7:0]    regVec_2854;
  reg        [7:0]    regVec_2855;
  reg        [7:0]    regVec_2856;
  reg        [7:0]    regVec_2857;
  reg        [7:0]    regVec_2858;
  reg        [7:0]    regVec_2859;
  reg        [7:0]    regVec_2860;
  reg        [7:0]    regVec_2861;
  reg        [7:0]    regVec_2862;
  reg        [7:0]    regVec_2863;
  reg        [7:0]    regVec_2864;
  reg        [7:0]    regVec_2865;
  reg        [7:0]    regVec_2866;
  reg        [7:0]    regVec_2867;
  reg        [7:0]    regVec_2868;
  reg        [7:0]    regVec_2869;
  reg        [7:0]    regVec_2870;
  reg        [7:0]    regVec_2871;
  reg        [7:0]    regVec_2872;
  reg        [7:0]    regVec_2873;
  reg        [7:0]    regVec_2874;
  reg        [7:0]    regVec_2875;
  reg        [7:0]    regVec_2876;
  reg        [7:0]    regVec_2877;
  reg        [7:0]    regVec_2878;
  reg        [7:0]    regVec_2879;
  reg        [7:0]    regVec_2880;
  reg        [7:0]    regVec_2881;
  reg        [7:0]    regVec_2882;
  reg        [7:0]    regVec_2883;
  reg        [7:0]    regVec_2884;
  reg        [7:0]    regVec_2885;
  reg        [7:0]    regVec_2886;
  reg        [7:0]    regVec_2887;
  reg        [7:0]    regVec_2888;
  reg        [7:0]    regVec_2889;
  reg        [7:0]    regVec_2890;
  reg        [7:0]    regVec_2891;
  reg        [7:0]    regVec_2892;
  reg        [7:0]    regVec_2893;
  reg        [7:0]    regVec_2894;
  reg        [7:0]    regVec_2895;
  reg        [7:0]    regVec_2896;
  reg        [7:0]    regVec_2897;
  reg        [7:0]    regVec_2898;
  reg        [7:0]    regVec_2899;
  reg        [7:0]    regVec_2900;
  reg        [7:0]    regVec_2901;
  reg        [7:0]    regVec_2902;
  reg        [7:0]    regVec_2903;
  reg        [7:0]    regVec_2904;
  reg        [7:0]    regVec_2905;
  reg        [7:0]    regVec_2906;
  reg        [7:0]    regVec_2907;
  reg        [7:0]    regVec_2908;
  reg        [7:0]    regVec_2909;
  reg        [7:0]    regVec_2910;
  reg        [7:0]    regVec_2911;
  reg        [7:0]    regVec_2912;
  reg        [7:0]    regVec_2913;
  reg        [7:0]    regVec_2914;
  reg        [7:0]    regVec_2915;
  reg        [7:0]    regVec_2916;
  reg        [7:0]    regVec_2917;
  reg        [7:0]    regVec_2918;
  reg        [7:0]    regVec_2919;
  reg        [7:0]    regVec_2920;
  reg        [7:0]    regVec_2921;
  reg        [7:0]    regVec_2922;
  reg        [7:0]    regVec_2923;
  reg        [7:0]    regVec_2924;
  reg        [7:0]    regVec_2925;
  reg        [7:0]    regVec_2926;
  reg        [7:0]    regVec_2927;
  reg        [7:0]    regVec_2928;
  reg        [7:0]    regVec_2929;
  reg        [7:0]    regVec_2930;
  reg        [7:0]    regVec_2931;
  reg        [7:0]    regVec_2932;
  reg        [7:0]    regVec_2933;
  reg        [7:0]    regVec_2934;
  reg        [7:0]    regVec_2935;
  reg        [7:0]    regVec_2936;
  reg        [7:0]    regVec_2937;
  reg        [7:0]    regVec_2938;
  reg        [7:0]    regVec_2939;
  reg        [7:0]    regVec_2940;
  reg        [7:0]    regVec_2941;
  reg        [7:0]    regVec_2942;
  reg        [7:0]    regVec_2943;
  reg        [7:0]    regVec_2944;
  reg        [7:0]    regVec_2945;
  reg        [7:0]    regVec_2946;
  reg        [7:0]    regVec_2947;
  reg        [7:0]    regVec_2948;
  reg        [7:0]    regVec_2949;
  reg        [7:0]    regVec_2950;
  reg        [7:0]    regVec_2951;
  reg        [7:0]    regVec_2952;
  reg        [7:0]    regVec_2953;
  reg        [7:0]    regVec_2954;
  reg        [7:0]    regVec_2955;
  reg        [7:0]    regVec_2956;
  reg        [7:0]    regVec_2957;
  reg        [7:0]    regVec_2958;
  reg        [7:0]    regVec_2959;
  reg        [7:0]    regVec_2960;
  reg        [7:0]    regVec_2961;
  reg        [7:0]    regVec_2962;
  reg        [7:0]    regVec_2963;
  reg        [7:0]    regVec_2964;
  reg        [7:0]    regVec_2965;
  reg        [7:0]    regVec_2966;
  reg        [7:0]    regVec_2967;
  reg        [7:0]    regVec_2968;
  reg        [7:0]    regVec_2969;
  reg        [7:0]    regVec_2970;
  reg        [7:0]    regVec_2971;
  reg        [7:0]    regVec_2972;
  reg        [7:0]    regVec_2973;
  reg        [7:0]    regVec_2974;
  reg        [7:0]    regVec_2975;
  reg        [7:0]    regVec_2976;
  reg        [7:0]    regVec_2977;
  reg        [7:0]    regVec_2978;
  reg        [7:0]    regVec_2979;
  reg        [7:0]    regVec_2980;
  reg        [7:0]    regVec_2981;
  reg        [7:0]    regVec_2982;
  reg        [7:0]    regVec_2983;
  reg        [7:0]    regVec_2984;
  reg        [7:0]    regVec_2985;
  reg        [7:0]    regVec_2986;
  reg        [7:0]    regVec_2987;
  reg        [7:0]    regVec_2988;
  reg        [7:0]    regVec_2989;
  reg        [7:0]    regVec_2990;
  reg        [7:0]    regVec_2991;
  reg        [7:0]    regVec_2992;
  reg        [7:0]    regVec_2993;
  reg        [7:0]    regVec_2994;
  reg        [7:0]    regVec_2995;
  reg        [7:0]    regVec_2996;
  reg        [7:0]    regVec_2997;
  reg        [7:0]    regVec_2998;
  reg        [7:0]    regVec_2999;
  reg        [7:0]    regVec_3000;
  reg        [7:0]    regVec_3001;
  reg        [7:0]    regVec_3002;
  reg        [7:0]    regVec_3003;
  reg        [7:0]    regVec_3004;
  reg        [7:0]    regVec_3005;
  reg        [7:0]    regVec_3006;
  reg        [7:0]    regVec_3007;
  reg        [7:0]    regVec_3008;
  reg        [7:0]    regVec_3009;
  reg        [7:0]    regVec_3010;
  reg        [7:0]    regVec_3011;
  reg        [7:0]    regVec_3012;
  reg        [7:0]    regVec_3013;
  reg        [7:0]    regVec_3014;
  reg        [7:0]    regVec_3015;
  reg        [7:0]    regVec_3016;
  reg        [7:0]    regVec_3017;
  reg        [7:0]    regVec_3018;
  reg        [7:0]    regVec_3019;
  reg        [7:0]    regVec_3020;
  reg        [7:0]    regVec_3021;
  reg        [7:0]    regVec_3022;
  reg        [7:0]    regVec_3023;
  reg        [7:0]    regVec_3024;
  reg        [7:0]    regVec_3025;
  reg        [7:0]    regVec_3026;
  reg        [7:0]    regVec_3027;
  reg        [7:0]    regVec_3028;
  reg        [7:0]    regVec_3029;
  reg        [7:0]    regVec_3030;
  reg        [7:0]    regVec_3031;
  reg        [7:0]    regVec_3032;
  reg        [7:0]    regVec_3033;
  reg        [7:0]    regVec_3034;
  reg        [7:0]    regVec_3035;
  reg        [7:0]    regVec_3036;
  reg        [7:0]    regVec_3037;
  reg        [7:0]    regVec_3038;
  reg        [7:0]    regVec_3039;
  reg        [7:0]    regVec_3040;
  reg        [7:0]    regVec_3041;
  reg        [7:0]    regVec_3042;
  reg        [7:0]    regVec_3043;
  reg        [7:0]    regVec_3044;
  reg        [7:0]    regVec_3045;
  reg        [7:0]    regVec_3046;
  reg        [7:0]    regVec_3047;
  reg        [7:0]    regVec_3048;
  reg        [7:0]    regVec_3049;
  reg        [7:0]    regVec_3050;
  reg        [7:0]    regVec_3051;
  reg        [7:0]    regVec_3052;
  reg        [7:0]    regVec_3053;
  reg        [7:0]    regVec_3054;
  reg        [7:0]    regVec_3055;
  reg        [7:0]    regVec_3056;
  reg        [7:0]    regVec_3057;
  reg        [7:0]    regVec_3058;
  reg        [7:0]    regVec_3059;
  reg        [7:0]    regVec_3060;
  reg        [7:0]    regVec_3061;
  reg        [7:0]    regVec_3062;
  reg        [7:0]    regVec_3063;
  reg        [7:0]    regVec_3064;
  reg        [7:0]    regVec_3065;
  reg        [7:0]    regVec_3066;
  reg        [7:0]    regVec_3067;
  reg        [7:0]    regVec_3068;
  reg        [7:0]    regVec_3069;
  reg        [7:0]    regVec_3070;
  reg        [7:0]    regVec_3071;
  reg        [7:0]    regVec_3072;
  reg        [7:0]    regVec_3073;
  reg        [7:0]    regVec_3074;
  reg        [7:0]    regVec_3075;
  reg        [7:0]    regVec_3076;
  reg        [7:0]    regVec_3077;
  reg        [7:0]    regVec_3078;
  reg        [7:0]    regVec_3079;
  reg        [7:0]    regVec_3080;
  reg        [7:0]    regVec_3081;
  reg        [7:0]    regVec_3082;
  reg        [7:0]    regVec_3083;
  reg        [7:0]    regVec_3084;
  reg        [7:0]    regVec_3085;
  reg        [7:0]    regVec_3086;
  reg        [7:0]    regVec_3087;
  reg        [7:0]    regVec_3088;
  reg        [7:0]    regVec_3089;
  reg        [7:0]    regVec_3090;
  reg        [7:0]    regVec_3091;
  reg        [7:0]    regVec_3092;
  reg        [7:0]    regVec_3093;
  reg        [7:0]    regVec_3094;
  reg        [7:0]    regVec_3095;
  reg        [7:0]    regVec_3096;
  reg        [7:0]    regVec_3097;
  reg        [7:0]    regVec_3098;
  reg        [7:0]    regVec_3099;
  reg        [7:0]    regVec_3100;
  reg        [7:0]    regVec_3101;
  reg        [7:0]    regVec_3102;
  reg        [7:0]    regVec_3103;
  reg        [7:0]    regVec_3104;
  reg        [7:0]    regVec_3105;
  reg        [7:0]    regVec_3106;
  reg        [7:0]    regVec_3107;
  reg        [7:0]    regVec_3108;
  reg        [7:0]    regVec_3109;
  reg        [7:0]    regVec_3110;
  reg        [7:0]    regVec_3111;
  reg        [7:0]    regVec_3112;
  reg        [7:0]    regVec_3113;
  reg        [7:0]    regVec_3114;
  reg        [7:0]    regVec_3115;
  reg        [7:0]    regVec_3116;
  reg        [7:0]    regVec_3117;
  reg        [7:0]    regVec_3118;
  reg        [7:0]    regVec_3119;
  reg        [7:0]    regVec_3120;
  reg        [7:0]    regVec_3121;
  reg        [7:0]    regVec_3122;
  reg        [7:0]    regVec_3123;
  reg        [7:0]    regVec_3124;
  reg        [7:0]    regVec_3125;
  reg        [7:0]    regVec_3126;
  reg        [7:0]    regVec_3127;
  reg        [7:0]    regVec_3128;
  reg        [7:0]    regVec_3129;
  reg        [7:0]    regVec_3130;
  reg        [7:0]    regVec_3131;
  reg        [7:0]    regVec_3132;
  reg        [7:0]    regVec_3133;
  reg        [7:0]    regVec_3134;
  reg        [7:0]    regVec_3135;
  reg        [7:0]    regVec_3136;
  reg        [7:0]    regVec_3137;
  reg        [7:0]    regVec_3138;
  reg        [7:0]    regVec_3139;
  reg        [7:0]    regVec_3140;
  reg        [7:0]    regVec_3141;
  reg        [7:0]    regVec_3142;
  reg        [7:0]    regVec_3143;
  reg        [7:0]    regVec_3144;
  reg        [7:0]    regVec_3145;
  reg        [7:0]    regVec_3146;
  reg        [7:0]    regVec_3147;
  reg        [7:0]    regVec_3148;
  reg        [7:0]    regVec_3149;
  reg        [7:0]    regVec_3150;
  reg        [7:0]    regVec_3151;
  reg        [7:0]    regVec_3152;
  reg        [7:0]    regVec_3153;
  reg        [7:0]    regVec_3154;
  reg        [7:0]    regVec_3155;
  reg        [7:0]    regVec_3156;
  reg        [7:0]    regVec_3157;
  reg        [7:0]    regVec_3158;
  reg        [7:0]    regVec_3159;
  reg        [7:0]    regVec_3160;
  reg        [7:0]    regVec_3161;
  reg        [7:0]    regVec_3162;
  reg        [7:0]    regVec_3163;
  reg        [7:0]    regVec_3164;
  reg        [7:0]    regVec_3165;
  reg        [7:0]    regVec_3166;
  reg        [7:0]    regVec_3167;
  reg        [7:0]    regVec_3168;
  reg        [7:0]    regVec_3169;
  reg        [7:0]    regVec_3170;
  reg        [7:0]    regVec_3171;
  reg        [7:0]    regVec_3172;
  reg        [7:0]    regVec_3173;
  reg        [7:0]    regVec_3174;
  reg        [7:0]    regVec_3175;
  reg        [7:0]    regVec_3176;
  reg        [7:0]    regVec_3177;
  reg        [7:0]    regVec_3178;
  reg        [7:0]    regVec_3179;
  reg        [7:0]    regVec_3180;
  reg        [7:0]    regVec_3181;
  reg        [7:0]    regVec_3182;
  reg        [7:0]    regVec_3183;
  reg        [7:0]    regVec_3184;
  reg        [7:0]    regVec_3185;
  reg        [7:0]    regVec_3186;
  reg        [7:0]    regVec_3187;
  reg        [7:0]    regVec_3188;
  reg        [7:0]    regVec_3189;
  reg        [7:0]    regVec_3190;
  reg        [7:0]    regVec_3191;
  reg        [7:0]    regVec_3192;
  reg        [7:0]    regVec_3193;
  reg        [7:0]    regVec_3194;
  reg        [7:0]    regVec_3195;
  reg        [7:0]    regVec_3196;
  reg        [7:0]    regVec_3197;
  reg        [7:0]    regVec_3198;
  reg        [7:0]    regVec_3199;
  reg        [7:0]    regVec_3200;
  reg        [7:0]    regVec_3201;
  reg        [7:0]    regVec_3202;
  reg        [7:0]    regVec_3203;
  reg        [7:0]    regVec_3204;
  reg        [7:0]    regVec_3205;
  reg        [7:0]    regVec_3206;
  reg        [7:0]    regVec_3207;
  reg        [7:0]    regVec_3208;
  reg        [7:0]    regVec_3209;
  reg        [7:0]    regVec_3210;
  reg        [7:0]    regVec_3211;
  reg        [7:0]    regVec_3212;
  reg        [7:0]    regVec_3213;
  reg        [7:0]    regVec_3214;
  reg        [7:0]    regVec_3215;
  reg        [7:0]    regVec_3216;
  reg        [7:0]    regVec_3217;
  reg        [7:0]    regVec_3218;
  reg        [7:0]    regVec_3219;
  reg        [7:0]    regVec_3220;
  reg        [7:0]    regVec_3221;
  reg        [7:0]    regVec_3222;
  reg        [7:0]    regVec_3223;
  reg        [7:0]    regVec_3224;
  reg        [7:0]    regVec_3225;
  reg        [7:0]    regVec_3226;
  reg        [7:0]    regVec_3227;
  reg        [7:0]    regVec_3228;
  reg        [7:0]    regVec_3229;
  reg        [7:0]    regVec_3230;
  reg        [7:0]    regVec_3231;
  reg        [7:0]    regVec_3232;
  reg        [7:0]    regVec_3233;
  reg        [7:0]    regVec_3234;
  reg        [7:0]    regVec_3235;
  reg        [7:0]    regVec_3236;
  reg        [7:0]    regVec_3237;
  reg        [7:0]    regVec_3238;
  reg        [7:0]    regVec_3239;
  reg        [7:0]    regVec_3240;
  reg        [7:0]    regVec_3241;
  reg        [7:0]    regVec_3242;
  reg        [7:0]    regVec_3243;
  reg        [7:0]    regVec_3244;
  reg        [7:0]    regVec_3245;
  reg        [7:0]    regVec_3246;
  reg        [7:0]    regVec_3247;
  reg        [7:0]    regVec_3248;
  reg        [7:0]    regVec_3249;
  reg        [7:0]    regVec_3250;
  reg        [7:0]    regVec_3251;
  reg        [7:0]    regVec_3252;
  reg        [7:0]    regVec_3253;
  reg        [7:0]    regVec_3254;
  reg        [7:0]    regVec_3255;
  reg        [7:0]    regVec_3256;
  reg        [7:0]    regVec_3257;
  reg        [7:0]    regVec_3258;
  reg        [7:0]    regVec_3259;
  reg        [7:0]    regVec_3260;
  reg        [7:0]    regVec_3261;
  reg        [7:0]    regVec_3262;
  reg        [7:0]    regVec_3263;
  reg        [7:0]    regVec_3264;
  reg        [7:0]    regVec_3265;
  reg        [7:0]    regVec_3266;
  reg        [7:0]    regVec_3267;
  reg        [7:0]    regVec_3268;
  reg        [7:0]    regVec_3269;
  reg        [7:0]    regVec_3270;
  reg        [7:0]    regVec_3271;
  reg        [7:0]    regVec_3272;
  reg        [7:0]    regVec_3273;
  reg        [7:0]    regVec_3274;
  reg        [7:0]    regVec_3275;
  reg        [7:0]    regVec_3276;
  reg        [7:0]    regVec_3277;
  reg        [7:0]    regVec_3278;
  reg        [7:0]    regVec_3279;
  reg        [7:0]    regVec_3280;
  reg        [7:0]    regVec_3281;
  reg        [7:0]    regVec_3282;
  reg        [7:0]    regVec_3283;
  reg        [7:0]    regVec_3284;
  reg        [7:0]    regVec_3285;
  reg        [7:0]    regVec_3286;
  reg        [7:0]    regVec_3287;
  reg        [7:0]    regVec_3288;
  reg        [7:0]    regVec_3289;
  reg        [7:0]    regVec_3290;
  reg        [7:0]    regVec_3291;
  reg        [7:0]    regVec_3292;
  reg        [7:0]    regVec_3293;
  reg        [7:0]    regVec_3294;
  reg        [7:0]    regVec_3295;
  reg        [7:0]    regVec_3296;
  reg        [7:0]    regVec_3297;
  reg        [7:0]    regVec_3298;
  reg        [7:0]    regVec_3299;
  reg        [7:0]    regVec_3300;
  reg        [7:0]    regVec_3301;
  reg        [7:0]    regVec_3302;
  reg        [7:0]    regVec_3303;
  reg        [7:0]    regVec_3304;
  reg        [7:0]    regVec_3305;
  reg        [7:0]    regVec_3306;
  reg        [7:0]    regVec_3307;
  reg        [7:0]    regVec_3308;
  reg        [7:0]    regVec_3309;
  reg        [7:0]    regVec_3310;
  reg        [7:0]    regVec_3311;
  reg        [7:0]    regVec_3312;
  reg        [7:0]    regVec_3313;
  reg        [7:0]    regVec_3314;
  reg        [7:0]    regVec_3315;
  reg        [7:0]    regVec_3316;
  reg        [7:0]    regVec_3317;
  reg        [7:0]    regVec_3318;
  reg        [7:0]    regVec_3319;
  reg        [7:0]    regVec_3320;
  reg        [7:0]    regVec_3321;
  reg        [7:0]    regVec_3322;
  reg        [7:0]    regVec_3323;
  reg        [7:0]    regVec_3324;
  reg        [7:0]    regVec_3325;
  reg        [7:0]    regVec_3326;
  reg        [7:0]    regVec_3327;
  reg        [7:0]    regVec_3328;
  reg        [7:0]    regVec_3329;
  reg        [7:0]    regVec_3330;
  reg        [7:0]    regVec_3331;
  reg        [7:0]    regVec_3332;
  reg        [7:0]    regVec_3333;
  reg        [7:0]    regVec_3334;
  reg        [7:0]    regVec_3335;
  reg        [7:0]    regVec_3336;
  reg        [7:0]    regVec_3337;
  reg        [7:0]    regVec_3338;
  reg        [7:0]    regVec_3339;
  reg        [7:0]    regVec_3340;
  reg        [7:0]    regVec_3341;
  reg        [7:0]    regVec_3342;
  reg        [7:0]    regVec_3343;
  reg        [7:0]    regVec_3344;
  reg        [7:0]    regVec_3345;
  reg        [7:0]    regVec_3346;
  reg        [7:0]    regVec_3347;
  reg        [7:0]    regVec_3348;
  reg        [7:0]    regVec_3349;
  reg        [7:0]    regVec_3350;
  reg        [7:0]    regVec_3351;
  reg        [7:0]    regVec_3352;
  reg        [7:0]    regVec_3353;
  reg        [7:0]    regVec_3354;
  reg        [7:0]    regVec_3355;
  reg        [7:0]    regVec_3356;
  reg        [7:0]    regVec_3357;
  reg        [7:0]    regVec_3358;
  reg        [7:0]    regVec_3359;
  reg        [7:0]    regVec_3360;
  reg        [7:0]    regVec_3361;
  reg        [7:0]    regVec_3362;
  reg        [7:0]    regVec_3363;
  reg        [7:0]    regVec_3364;
  reg        [7:0]    regVec_3365;
  reg        [7:0]    regVec_3366;
  reg        [7:0]    regVec_3367;
  reg        [7:0]    regVec_3368;
  reg        [7:0]    regVec_3369;
  reg        [7:0]    regVec_3370;
  reg        [7:0]    regVec_3371;
  reg        [7:0]    regVec_3372;
  reg        [7:0]    regVec_3373;
  reg        [7:0]    regVec_3374;
  reg        [7:0]    regVec_3375;
  reg        [7:0]    regVec_3376;
  reg        [7:0]    regVec_3377;
  reg        [7:0]    regVec_3378;
  reg        [7:0]    regVec_3379;
  reg        [7:0]    regVec_3380;
  reg        [7:0]    regVec_3381;
  reg        [7:0]    regVec_3382;
  reg        [7:0]    regVec_3383;
  reg        [7:0]    regVec_3384;
  reg        [7:0]    regVec_3385;
  reg        [7:0]    regVec_3386;
  reg        [7:0]    regVec_3387;
  reg        [7:0]    regVec_3388;
  reg        [7:0]    regVec_3389;
  reg        [7:0]    regVec_3390;
  reg        [7:0]    regVec_3391;
  reg        [7:0]    regVec_3392;
  reg        [7:0]    regVec_3393;
  reg        [7:0]    regVec_3394;
  reg        [7:0]    regVec_3395;
  reg        [7:0]    regVec_3396;
  reg        [7:0]    regVec_3397;
  reg        [7:0]    regVec_3398;
  reg        [7:0]    regVec_3399;
  reg        [7:0]    regVec_3400;
  reg        [7:0]    regVec_3401;
  reg        [7:0]    regVec_3402;
  reg        [7:0]    regVec_3403;
  reg        [7:0]    regVec_3404;
  reg        [7:0]    regVec_3405;
  reg        [7:0]    regVec_3406;
  reg        [7:0]    regVec_3407;
  reg        [7:0]    regVec_3408;
  reg        [7:0]    regVec_3409;
  reg        [7:0]    regVec_3410;
  reg        [7:0]    regVec_3411;
  reg        [7:0]    regVec_3412;
  reg        [7:0]    regVec_3413;
  reg        [7:0]    regVec_3414;
  reg        [7:0]    regVec_3415;
  reg        [7:0]    regVec_3416;
  reg        [7:0]    regVec_3417;
  reg        [7:0]    regVec_3418;
  reg        [7:0]    regVec_3419;
  reg        [7:0]    regVec_3420;
  reg        [7:0]    regVec_3421;
  reg        [7:0]    regVec_3422;
  reg        [7:0]    regVec_3423;
  reg        [7:0]    regVec_3424;
  reg        [7:0]    regVec_3425;
  reg        [7:0]    regVec_3426;
  reg        [7:0]    regVec_3427;
  reg        [7:0]    regVec_3428;
  reg        [7:0]    regVec_3429;
  reg        [7:0]    regVec_3430;
  reg        [7:0]    regVec_3431;
  reg        [7:0]    regVec_3432;
  reg        [7:0]    regVec_3433;
  reg        [7:0]    regVec_3434;
  reg        [7:0]    regVec_3435;
  reg        [7:0]    regVec_3436;
  reg        [7:0]    regVec_3437;
  reg        [7:0]    regVec_3438;
  reg        [7:0]    regVec_3439;
  reg        [7:0]    regVec_3440;
  reg        [7:0]    regVec_3441;
  reg        [7:0]    regVec_3442;
  reg        [7:0]    regVec_3443;
  reg        [7:0]    regVec_3444;
  reg        [7:0]    regVec_3445;
  reg        [7:0]    regVec_3446;
  reg        [7:0]    regVec_3447;
  reg        [7:0]    regVec_3448;
  reg        [7:0]    regVec_3449;
  reg        [7:0]    regVec_3450;
  reg        [7:0]    regVec_3451;
  reg        [7:0]    regVec_3452;
  reg        [7:0]    regVec_3453;
  reg        [7:0]    regVec_3454;
  reg        [7:0]    regVec_3455;
  reg        [7:0]    regVec_3456;
  reg        [7:0]    regVec_3457;
  reg        [7:0]    regVec_3458;
  reg        [7:0]    regVec_3459;
  reg        [7:0]    regVec_3460;
  reg        [7:0]    regVec_3461;
  reg        [7:0]    regVec_3462;
  reg        [7:0]    regVec_3463;
  reg        [7:0]    regVec_3464;
  reg        [7:0]    regVec_3465;
  reg        [7:0]    regVec_3466;
  reg        [7:0]    regVec_3467;
  reg        [7:0]    regVec_3468;
  reg        [7:0]    regVec_3469;
  reg        [7:0]    regVec_3470;
  reg        [7:0]    regVec_3471;
  reg        [7:0]    regVec_3472;
  reg        [7:0]    regVec_3473;
  reg        [7:0]    regVec_3474;
  reg        [7:0]    regVec_3475;
  reg        [7:0]    regVec_3476;
  reg        [7:0]    regVec_3477;
  reg        [7:0]    regVec_3478;
  reg        [7:0]    regVec_3479;
  reg        [7:0]    regVec_3480;
  reg        [7:0]    regVec_3481;
  reg        [7:0]    regVec_3482;
  reg        [7:0]    regVec_3483;
  reg        [7:0]    regVec_3484;
  reg        [7:0]    regVec_3485;
  reg        [7:0]    regVec_3486;
  reg        [7:0]    regVec_3487;
  reg        [7:0]    regVec_3488;
  reg        [7:0]    regVec_3489;
  reg        [7:0]    regVec_3490;
  reg        [7:0]    regVec_3491;
  reg        [7:0]    regVec_3492;
  reg        [7:0]    regVec_3493;
  reg        [7:0]    regVec_3494;
  reg        [7:0]    regVec_3495;
  reg        [7:0]    regVec_3496;
  reg        [7:0]    regVec_3497;
  reg        [7:0]    regVec_3498;
  reg        [7:0]    regVec_3499;
  reg        [7:0]    regVec_3500;
  reg        [7:0]    regVec_3501;
  reg        [7:0]    regVec_3502;
  reg        [7:0]    regVec_3503;
  reg        [7:0]    regVec_3504;
  reg        [7:0]    regVec_3505;
  reg        [7:0]    regVec_3506;
  reg        [7:0]    regVec_3507;
  reg        [7:0]    regVec_3508;
  reg        [7:0]    regVec_3509;
  reg        [7:0]    regVec_3510;
  reg        [7:0]    regVec_3511;
  reg        [7:0]    regVec_3512;
  reg        [7:0]    regVec_3513;
  reg        [7:0]    regVec_3514;
  reg        [7:0]    regVec_3515;
  reg        [7:0]    regVec_3516;
  reg        [7:0]    regVec_3517;
  reg        [7:0]    regVec_3518;
  reg        [7:0]    regVec_3519;
  reg        [7:0]    regVec_3520;
  reg        [7:0]    regVec_3521;
  reg        [7:0]    regVec_3522;
  reg        [7:0]    regVec_3523;
  reg        [7:0]    regVec_3524;
  reg        [7:0]    regVec_3525;
  reg        [7:0]    regVec_3526;
  reg        [7:0]    regVec_3527;
  reg        [7:0]    regVec_3528;
  reg        [7:0]    regVec_3529;
  reg        [7:0]    regVec_3530;
  reg        [7:0]    regVec_3531;
  reg        [7:0]    regVec_3532;
  reg        [7:0]    regVec_3533;
  reg        [7:0]    regVec_3534;
  reg        [7:0]    regVec_3535;
  reg        [7:0]    regVec_3536;
  reg        [7:0]    regVec_3537;
  reg        [7:0]    regVec_3538;
  reg        [7:0]    regVec_3539;
  reg        [7:0]    regVec_3540;
  reg        [7:0]    regVec_3541;
  reg        [7:0]    regVec_3542;
  reg        [7:0]    regVec_3543;
  reg        [7:0]    regVec_3544;
  reg        [7:0]    regVec_3545;
  reg        [7:0]    regVec_3546;
  reg        [7:0]    regVec_3547;
  reg        [7:0]    regVec_3548;
  reg        [7:0]    regVec_3549;
  reg        [7:0]    regVec_3550;
  reg        [7:0]    regVec_3551;
  reg        [7:0]    regVec_3552;
  reg        [7:0]    regVec_3553;
  reg        [7:0]    regVec_3554;
  reg        [7:0]    regVec_3555;
  reg        [7:0]    regVec_3556;
  reg        [7:0]    regVec_3557;
  reg        [7:0]    regVec_3558;
  reg        [7:0]    regVec_3559;
  reg        [7:0]    regVec_3560;
  reg        [7:0]    regVec_3561;
  reg        [7:0]    regVec_3562;
  reg        [7:0]    regVec_3563;
  reg        [7:0]    regVec_3564;
  reg        [7:0]    regVec_3565;
  reg        [7:0]    regVec_3566;
  reg        [7:0]    regVec_3567;
  reg        [7:0]    regVec_3568;
  reg        [7:0]    regVec_3569;
  reg        [7:0]    regVec_3570;
  reg        [7:0]    regVec_3571;
  reg        [7:0]    regVec_3572;
  reg        [7:0]    regVec_3573;
  reg        [7:0]    regVec_3574;
  reg        [7:0]    regVec_3575;
  reg        [7:0]    regVec_3576;
  reg        [7:0]    regVec_3577;
  reg        [7:0]    regVec_3578;
  reg        [7:0]    regVec_3579;
  reg        [7:0]    regVec_3580;
  reg        [7:0]    regVec_3581;
  reg        [7:0]    regVec_3582;
  reg        [7:0]    regVec_3583;
  reg        [7:0]    regVec_3584;
  reg        [7:0]    regVec_3585;
  reg        [7:0]    regVec_3586;
  reg        [7:0]    regVec_3587;
  reg        [7:0]    regVec_3588;
  reg        [7:0]    regVec_3589;
  reg        [7:0]    regVec_3590;
  reg        [7:0]    regVec_3591;
  reg        [7:0]    regVec_3592;
  reg        [7:0]    regVec_3593;
  reg        [7:0]    regVec_3594;
  reg        [7:0]    regVec_3595;
  reg        [7:0]    regVec_3596;
  reg        [7:0]    regVec_3597;
  reg        [7:0]    regVec_3598;
  reg        [7:0]    regVec_3599;
  reg        [7:0]    regVec_3600;
  reg        [7:0]    regVec_3601;
  reg        [7:0]    regVec_3602;
  reg        [7:0]    regVec_3603;
  reg        [7:0]    regVec_3604;
  reg        [7:0]    regVec_3605;
  reg        [7:0]    regVec_3606;
  reg        [7:0]    regVec_3607;
  reg        [7:0]    regVec_3608;
  reg        [7:0]    regVec_3609;
  reg        [7:0]    regVec_3610;
  reg        [7:0]    regVec_3611;
  reg        [7:0]    regVec_3612;
  reg        [7:0]    regVec_3613;
  reg        [7:0]    regVec_3614;
  reg        [7:0]    regVec_3615;
  reg        [7:0]    regVec_3616;
  reg        [7:0]    regVec_3617;
  reg        [7:0]    regVec_3618;
  reg        [7:0]    regVec_3619;
  reg        [7:0]    regVec_3620;
  reg        [7:0]    regVec_3621;
  reg        [7:0]    regVec_3622;
  reg        [7:0]    regVec_3623;
  reg        [7:0]    regVec_3624;
  reg        [7:0]    regVec_3625;
  reg        [7:0]    regVec_3626;
  reg        [7:0]    regVec_3627;
  reg        [7:0]    regVec_3628;
  reg        [7:0]    regVec_3629;
  reg        [7:0]    regVec_3630;
  reg        [7:0]    regVec_3631;
  reg        [7:0]    regVec_3632;
  reg        [7:0]    regVec_3633;
  reg        [7:0]    regVec_3634;
  reg        [7:0]    regVec_3635;
  reg        [7:0]    regVec_3636;
  reg        [7:0]    regVec_3637;
  reg        [7:0]    regVec_3638;
  reg        [7:0]    regVec_3639;
  reg        [7:0]    regVec_3640;
  reg        [7:0]    regVec_3641;
  reg        [7:0]    regVec_3642;
  reg        [7:0]    regVec_3643;
  reg        [7:0]    regVec_3644;
  reg        [7:0]    regVec_3645;
  reg        [7:0]    regVec_3646;
  reg        [7:0]    regVec_3647;
  reg        [7:0]    regVec_3648;
  reg        [7:0]    regVec_3649;
  reg        [7:0]    regVec_3650;
  reg        [7:0]    regVec_3651;
  reg        [7:0]    regVec_3652;
  reg        [7:0]    regVec_3653;
  reg        [7:0]    regVec_3654;
  reg        [7:0]    regVec_3655;
  reg        [7:0]    regVec_3656;
  reg        [7:0]    regVec_3657;
  reg        [7:0]    regVec_3658;
  reg        [7:0]    regVec_3659;
  reg        [7:0]    regVec_3660;
  reg        [7:0]    regVec_3661;
  reg        [7:0]    regVec_3662;
  reg        [7:0]    regVec_3663;
  reg        [7:0]    regVec_3664;
  reg        [7:0]    regVec_3665;
  reg        [7:0]    regVec_3666;
  reg        [7:0]    regVec_3667;
  reg        [7:0]    regVec_3668;
  reg        [7:0]    regVec_3669;
  reg        [7:0]    regVec_3670;
  reg        [7:0]    regVec_3671;
  reg        [7:0]    regVec_3672;
  reg        [7:0]    regVec_3673;
  reg        [7:0]    regVec_3674;
  reg        [7:0]    regVec_3675;
  reg        [7:0]    regVec_3676;
  reg        [7:0]    regVec_3677;
  reg        [7:0]    regVec_3678;
  reg        [7:0]    regVec_3679;
  reg        [7:0]    regVec_3680;
  reg        [7:0]    regVec_3681;
  reg        [7:0]    regVec_3682;
  reg        [7:0]    regVec_3683;
  reg        [7:0]    regVec_3684;
  reg        [7:0]    regVec_3685;
  reg        [7:0]    regVec_3686;
  reg        [7:0]    regVec_3687;
  reg        [7:0]    regVec_3688;
  reg        [7:0]    regVec_3689;
  reg        [7:0]    regVec_3690;
  reg        [7:0]    regVec_3691;
  reg        [7:0]    regVec_3692;
  reg        [7:0]    regVec_3693;
  reg        [7:0]    regVec_3694;
  reg        [7:0]    regVec_3695;
  reg        [7:0]    regVec_3696;
  reg        [7:0]    regVec_3697;
  reg        [7:0]    regVec_3698;
  reg        [7:0]    regVec_3699;
  reg        [7:0]    regVec_3700;
  reg        [7:0]    regVec_3701;
  reg        [7:0]    regVec_3702;
  reg        [7:0]    regVec_3703;
  reg        [7:0]    regVec_3704;
  reg        [7:0]    regVec_3705;
  reg        [7:0]    regVec_3706;
  reg        [7:0]    regVec_3707;
  reg        [7:0]    regVec_3708;
  reg        [7:0]    regVec_3709;
  reg        [7:0]    regVec_3710;
  reg        [7:0]    regVec_3711;
  reg        [7:0]    regVec_3712;
  reg        [7:0]    regVec_3713;
  reg        [7:0]    regVec_3714;
  reg        [7:0]    regVec_3715;
  reg        [7:0]    regVec_3716;
  reg        [7:0]    regVec_3717;
  reg        [7:0]    regVec_3718;
  reg        [7:0]    regVec_3719;
  reg        [7:0]    regVec_3720;
  reg        [7:0]    regVec_3721;
  reg        [7:0]    regVec_3722;
  reg        [7:0]    regVec_3723;
  reg        [7:0]    regVec_3724;
  reg        [7:0]    regVec_3725;
  reg        [7:0]    regVec_3726;
  reg        [7:0]    regVec_3727;
  reg        [7:0]    regVec_3728;
  reg        [7:0]    regVec_3729;
  reg        [7:0]    regVec_3730;
  reg        [7:0]    regVec_3731;
  reg        [7:0]    regVec_3732;
  reg        [7:0]    regVec_3733;
  reg        [7:0]    regVec_3734;
  reg        [7:0]    regVec_3735;
  reg        [7:0]    regVec_3736;
  reg        [7:0]    regVec_3737;
  reg        [7:0]    regVec_3738;
  reg        [7:0]    regVec_3739;
  reg        [7:0]    regVec_3740;
  reg        [7:0]    regVec_3741;
  reg        [7:0]    regVec_3742;
  reg        [7:0]    regVec_3743;
  reg        [7:0]    regVec_3744;
  reg        [7:0]    regVec_3745;
  reg        [7:0]    regVec_3746;
  reg        [7:0]    regVec_3747;
  reg        [7:0]    regVec_3748;
  reg        [7:0]    regVec_3749;
  reg        [7:0]    regVec_3750;
  reg        [7:0]    regVec_3751;
  reg        [7:0]    regVec_3752;
  reg        [7:0]    regVec_3753;
  reg        [7:0]    regVec_3754;
  reg        [7:0]    regVec_3755;
  reg        [7:0]    regVec_3756;
  reg        [7:0]    regVec_3757;
  reg        [7:0]    regVec_3758;
  reg        [7:0]    regVec_3759;
  reg        [7:0]    regVec_3760;
  reg        [7:0]    regVec_3761;
  reg        [7:0]    regVec_3762;
  reg        [7:0]    regVec_3763;
  reg        [7:0]    regVec_3764;
  reg        [7:0]    regVec_3765;
  reg        [7:0]    regVec_3766;
  reg        [7:0]    regVec_3767;
  reg        [7:0]    regVec_3768;
  reg        [7:0]    regVec_3769;
  reg        [7:0]    regVec_3770;
  reg        [7:0]    regVec_3771;
  reg        [7:0]    regVec_3772;
  reg        [7:0]    regVec_3773;
  reg        [7:0]    regVec_3774;
  reg        [7:0]    regVec_3775;
  reg        [7:0]    regVec_3776;
  reg        [7:0]    regVec_3777;
  reg        [7:0]    regVec_3778;
  reg        [7:0]    regVec_3779;
  reg        [7:0]    regVec_3780;
  reg        [7:0]    regVec_3781;
  reg        [7:0]    regVec_3782;
  reg        [7:0]    regVec_3783;
  reg        [7:0]    regVec_3784;
  reg        [7:0]    regVec_3785;
  reg        [7:0]    regVec_3786;
  reg        [7:0]    regVec_3787;
  reg        [7:0]    regVec_3788;
  reg        [7:0]    regVec_3789;
  reg        [7:0]    regVec_3790;
  reg        [7:0]    regVec_3791;
  reg        [7:0]    regVec_3792;
  reg        [7:0]    regVec_3793;
  reg        [7:0]    regVec_3794;
  reg        [7:0]    regVec_3795;
  reg        [7:0]    regVec_3796;
  reg        [7:0]    regVec_3797;
  reg        [7:0]    regVec_3798;
  reg        [7:0]    regVec_3799;
  reg        [7:0]    regVec_3800;
  reg        [7:0]    regVec_3801;
  reg        [7:0]    regVec_3802;
  reg        [7:0]    regVec_3803;
  reg        [7:0]    regVec_3804;
  reg        [7:0]    regVec_3805;
  reg        [7:0]    regVec_3806;
  reg        [7:0]    regVec_3807;
  reg        [7:0]    regVec_3808;
  reg        [7:0]    regVec_3809;
  reg        [7:0]    regVec_3810;
  reg        [7:0]    regVec_3811;
  reg        [7:0]    regVec_3812;
  reg        [7:0]    regVec_3813;
  reg        [7:0]    regVec_3814;
  reg        [7:0]    regVec_3815;
  reg        [7:0]    regVec_3816;
  reg        [7:0]    regVec_3817;
  reg        [7:0]    regVec_3818;
  reg        [7:0]    regVec_3819;
  reg        [7:0]    regVec_3820;
  reg        [7:0]    regVec_3821;
  reg        [7:0]    regVec_3822;
  reg        [7:0]    regVec_3823;
  reg        [7:0]    regVec_3824;
  reg        [7:0]    regVec_3825;
  reg        [7:0]    regVec_3826;
  reg        [7:0]    regVec_3827;
  reg        [7:0]    regVec_3828;
  reg        [7:0]    regVec_3829;
  reg        [7:0]    regVec_3830;
  reg        [7:0]    regVec_3831;
  reg        [7:0]    regVec_3832;
  reg        [7:0]    regVec_3833;
  reg        [7:0]    regVec_3834;
  reg        [7:0]    regVec_3835;
  reg        [7:0]    regVec_3836;
  reg        [7:0]    regVec_3837;
  reg        [7:0]    regVec_3838;
  reg        [7:0]    regVec_3839;
  reg        [7:0]    regVec_3840;
  reg        [7:0]    regVec_3841;
  reg        [7:0]    regVec_3842;
  reg        [7:0]    regVec_3843;
  reg        [7:0]    regVec_3844;
  reg        [7:0]    regVec_3845;
  reg        [7:0]    regVec_3846;
  reg        [7:0]    regVec_3847;
  reg        [7:0]    regVec_3848;
  reg        [7:0]    regVec_3849;
  reg        [7:0]    regVec_3850;
  reg        [7:0]    regVec_3851;
  reg        [7:0]    regVec_3852;
  reg        [7:0]    regVec_3853;
  reg        [7:0]    regVec_3854;
  reg        [7:0]    regVec_3855;
  reg        [7:0]    regVec_3856;
  reg        [7:0]    regVec_3857;
  reg        [7:0]    regVec_3858;
  reg        [7:0]    regVec_3859;
  reg        [7:0]    regVec_3860;
  reg        [7:0]    regVec_3861;
  reg        [7:0]    regVec_3862;
  reg        [7:0]    regVec_3863;
  reg        [7:0]    regVec_3864;
  reg        [7:0]    regVec_3865;
  reg        [7:0]    regVec_3866;
  reg        [7:0]    regVec_3867;
  reg        [7:0]    regVec_3868;
  reg        [7:0]    regVec_3869;
  reg        [7:0]    regVec_3870;
  reg        [7:0]    regVec_3871;
  reg        [7:0]    regVec_3872;
  reg        [7:0]    regVec_3873;
  reg        [7:0]    regVec_3874;
  reg        [7:0]    regVec_3875;
  reg        [7:0]    regVec_3876;
  reg        [7:0]    regVec_3877;
  reg        [7:0]    regVec_3878;
  reg        [7:0]    regVec_3879;
  reg        [7:0]    regVec_3880;
  reg        [7:0]    regVec_3881;
  reg        [7:0]    regVec_3882;
  reg        [7:0]    regVec_3883;
  reg        [7:0]    regVec_3884;
  reg        [7:0]    regVec_3885;
  reg        [7:0]    regVec_3886;
  reg        [7:0]    regVec_3887;
  reg        [7:0]    regVec_3888;
  reg        [7:0]    regVec_3889;
  reg        [7:0]    regVec_3890;
  reg        [7:0]    regVec_3891;
  reg        [7:0]    regVec_3892;
  reg        [7:0]    regVec_3893;
  reg        [7:0]    regVec_3894;
  reg        [7:0]    regVec_3895;
  reg        [7:0]    regVec_3896;
  reg        [7:0]    regVec_3897;
  reg        [7:0]    regVec_3898;
  reg        [7:0]    regVec_3899;
  reg        [7:0]    regVec_3900;
  reg        [7:0]    regVec_3901;
  reg        [7:0]    regVec_3902;
  reg        [7:0]    regVec_3903;
  reg        [7:0]    regVec_3904;
  reg        [7:0]    regVec_3905;
  reg        [7:0]    regVec_3906;
  reg        [7:0]    regVec_3907;
  reg        [7:0]    regVec_3908;
  reg        [7:0]    regVec_3909;
  reg        [7:0]    regVec_3910;
  reg        [7:0]    regVec_3911;
  reg        [7:0]    regVec_3912;
  reg        [7:0]    regVec_3913;
  reg        [7:0]    regVec_3914;
  reg        [7:0]    regVec_3915;
  reg        [7:0]    regVec_3916;
  reg        [7:0]    regVec_3917;
  reg        [7:0]    regVec_3918;
  reg        [7:0]    regVec_3919;
  reg        [7:0]    regVec_3920;
  reg        [7:0]    regVec_3921;
  reg        [7:0]    regVec_3922;
  reg        [7:0]    regVec_3923;
  reg        [7:0]    regVec_3924;
  reg        [7:0]    regVec_3925;
  reg        [7:0]    regVec_3926;
  reg        [7:0]    regVec_3927;
  reg        [7:0]    regVec_3928;
  reg        [7:0]    regVec_3929;
  reg        [7:0]    regVec_3930;
  reg        [7:0]    regVec_3931;
  reg        [7:0]    regVec_3932;
  reg        [7:0]    regVec_3933;
  reg        [7:0]    regVec_3934;
  reg        [7:0]    regVec_3935;
  reg        [7:0]    regVec_3936;
  reg        [7:0]    regVec_3937;
  reg        [7:0]    regVec_3938;
  reg        [7:0]    regVec_3939;
  reg        [7:0]    regVec_3940;
  reg        [7:0]    regVec_3941;
  reg        [7:0]    regVec_3942;
  reg        [7:0]    regVec_3943;
  reg        [7:0]    regVec_3944;
  reg        [7:0]    regVec_3945;
  reg        [7:0]    regVec_3946;
  reg        [7:0]    regVec_3947;
  reg        [7:0]    regVec_3948;
  reg        [7:0]    regVec_3949;
  reg        [7:0]    regVec_3950;
  reg        [7:0]    regVec_3951;
  reg        [7:0]    regVec_3952;
  reg        [7:0]    regVec_3953;
  reg        [7:0]    regVec_3954;
  reg        [7:0]    regVec_3955;
  reg        [7:0]    regVec_3956;
  reg        [7:0]    regVec_3957;
  reg        [7:0]    regVec_3958;
  reg        [7:0]    regVec_3959;
  reg        [7:0]    regVec_3960;
  reg        [7:0]    regVec_3961;
  reg        [7:0]    regVec_3962;
  reg        [7:0]    regVec_3963;
  reg        [7:0]    regVec_3964;
  reg        [7:0]    regVec_3965;
  reg        [7:0]    regVec_3966;
  reg        [7:0]    regVec_3967;
  reg        [7:0]    regVec_3968;
  reg        [7:0]    regVec_3969;
  reg        [7:0]    regVec_3970;
  reg        [7:0]    regVec_3971;
  reg        [7:0]    regVec_3972;
  reg        [7:0]    regVec_3973;
  reg        [7:0]    regVec_3974;
  reg        [7:0]    regVec_3975;
  reg        [7:0]    regVec_3976;
  reg        [7:0]    regVec_3977;
  reg        [7:0]    regVec_3978;
  reg        [7:0]    regVec_3979;
  reg        [7:0]    regVec_3980;
  reg        [7:0]    regVec_3981;
  reg        [7:0]    regVec_3982;
  reg        [7:0]    regVec_3983;
  reg        [7:0]    regVec_3984;
  reg        [7:0]    regVec_3985;
  reg        [7:0]    regVec_3986;
  reg        [7:0]    regVec_3987;
  reg        [7:0]    regVec_3988;
  reg        [7:0]    regVec_3989;
  reg        [7:0]    regVec_3990;
  reg        [7:0]    regVec_3991;
  reg        [7:0]    regVec_3992;
  reg        [7:0]    regVec_3993;
  reg        [7:0]    regVec_3994;
  reg        [7:0]    regVec_3995;
  reg        [7:0]    regVec_3996;
  reg        [7:0]    regVec_3997;
  reg        [7:0]    regVec_3998;
  reg        [7:0]    regVec_3999;
  reg        [7:0]    regVec_4000;
  reg        [7:0]    regVec_4001;
  reg        [7:0]    regVec_4002;
  reg        [7:0]    regVec_4003;
  reg        [7:0]    regVec_4004;
  reg        [7:0]    regVec_4005;
  reg        [7:0]    regVec_4006;
  reg        [7:0]    regVec_4007;
  reg        [7:0]    regVec_4008;
  reg        [7:0]    regVec_4009;
  reg        [7:0]    regVec_4010;
  reg        [7:0]    regVec_4011;
  reg        [7:0]    regVec_4012;
  reg        [7:0]    regVec_4013;
  reg        [7:0]    regVec_4014;
  reg        [7:0]    regVec_4015;
  reg        [7:0]    regVec_4016;
  reg        [7:0]    regVec_4017;
  reg        [7:0]    regVec_4018;
  reg        [7:0]    regVec_4019;
  reg        [7:0]    regVec_4020;
  reg        [7:0]    regVec_4021;
  reg        [7:0]    regVec_4022;
  reg        [7:0]    regVec_4023;
  reg        [7:0]    regVec_4024;
  reg        [7:0]    regVec_4025;
  reg        [7:0]    regVec_4026;
  reg        [7:0]    regVec_4027;
  reg        [7:0]    regVec_4028;
  reg        [7:0]    regVec_4029;
  reg        [7:0]    regVec_4030;
  reg        [7:0]    regVec_4031;
  reg        [7:0]    regVec_4032;
  reg        [7:0]    regVec_4033;
  reg        [7:0]    regVec_4034;
  reg        [7:0]    regVec_4035;
  reg        [7:0]    regVec_4036;
  reg        [7:0]    regVec_4037;
  reg        [7:0]    regVec_4038;
  reg        [7:0]    regVec_4039;
  reg        [7:0]    regVec_4040;
  reg        [7:0]    regVec_4041;
  reg        [7:0]    regVec_4042;
  reg        [7:0]    regVec_4043;
  reg        [7:0]    regVec_4044;
  reg        [7:0]    regVec_4045;
  reg        [7:0]    regVec_4046;
  reg        [7:0]    regVec_4047;
  reg        [7:0]    regVec_4048;
  reg        [7:0]    regVec_4049;
  reg        [7:0]    regVec_4050;
  reg        [7:0]    regVec_4051;
  reg        [7:0]    regVec_4052;
  reg        [7:0]    regVec_4053;
  reg        [7:0]    regVec_4054;
  reg        [7:0]    regVec_4055;
  reg        [7:0]    regVec_4056;
  reg        [7:0]    regVec_4057;
  reg        [7:0]    regVec_4058;
  reg        [7:0]    regVec_4059;
  reg        [7:0]    regVec_4060;
  reg        [7:0]    regVec_4061;
  reg        [7:0]    regVec_4062;
  reg        [7:0]    regVec_4063;
  reg        [7:0]    regVec_4064;
  reg        [7:0]    regVec_4065;
  reg        [7:0]    regVec_4066;
  reg        [7:0]    regVec_4067;
  reg        [7:0]    regVec_4068;
  reg        [7:0]    regVec_4069;
  reg        [7:0]    regVec_4070;
  reg        [7:0]    regVec_4071;
  reg        [7:0]    regVec_4072;
  reg        [7:0]    regVec_4073;
  reg        [7:0]    regVec_4074;
  reg        [7:0]    regVec_4075;
  reg        [7:0]    regVec_4076;
  reg        [7:0]    regVec_4077;
  reg        [7:0]    regVec_4078;
  reg        [7:0]    regVec_4079;
  reg        [7:0]    regVec_4080;
  reg        [7:0]    regVec_4081;
  reg        [7:0]    regVec_4082;
  reg        [7:0]    regVec_4083;
  reg        [7:0]    regVec_4084;
  reg        [7:0]    regVec_4085;
  reg        [7:0]    regVec_4086;
  reg        [7:0]    regVec_4087;
  reg        [7:0]    regVec_4088;
  reg        [7:0]    regVec_4089;
  reg        [7:0]    regVec_4090;
  reg        [7:0]    regVec_4091;
  reg        [7:0]    regVec_4092;
  reg        [7:0]    regVec_4093;
  reg        [7:0]    regVec_4094;
  reg        [7:0]    regVec_4095;
  reg        [11:0]   regAwAddr /* verilator public */ ;
  reg        [3:0]    regAwId;
  reg        [3:0]    regAwRegion;
  reg        [7:0]    regAwLen;
  reg        [2:0]    regAwSize;
  reg        [1:0]    regAwBrust;
  reg        [0:0]    regAwLock;
  reg        [3:0]    regAwCache;
  reg        [3:0]    regAwQos;
  reg        [0:0]    regAwUser;
  reg        [2:0]    regAwProt;
  reg        [11:0]   regArAddr;
  reg        [3:0]    regArId;
  reg        [3:0]    regArRegion;
  reg        [7:0]    regArLen;
  reg        [2:0]    regArSize;
  reg        [1:0]    regArBrust;
  reg        [0:0]    regArLock;
  reg        [3:0]    regArCache;
  reg        [3:0]    regArQos;
  reg        [0:0]    regArUser;
  reg        [2:0]    regArProt;
  reg                 updataAw;
  reg                 writeSuccess;
  reg                 updataAr;
  reg                 rFireCounter_willIncrement;
  wire                rFireCounter_willClear;
  reg        [12:0]   rFireCounter_valueNext;
  reg        [12:0]   rFireCounter_value;
  wire                rFireCounter_willOverflowIfInc;
  wire                rFireCounter_willOverflow;
  wire       [0:0]    bytePerWord;
  reg                 AwArConflict;
  wire                resetSignalValue;
  wire                when_Axi4_transmission_l66;
  wire                when_Axi4_transmission_l68;
  wire                when_Axi4_transmission_l72;
  wire                when_Axi4_transmission_l91;
  wire                when_Axi4_transmission_l92;
  wire       [4095:0] _zz_1;
  wire       [7:0]    _zz_regVec_0;
  wire       [4095:0] _zz_2;
  wire       [7:0]    _zz_regVec_0_1;
  reg        [11:0]   Axi4Incr_result;
  wire       [0:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [1:0]    Axi4Incr_wrapCase;
  wire                when_Axi4_transmission_l128;
  wire                when_Axi4_transmission_l132;
  wire                when_Axi4_transmission_l138;
  wire                when_Axi4_transmission_l140;
  wire                when_Axi4_transmission_l144;
  wire                when_Axi4_transmission_l171;
  reg        [11:0]   Axi4Incr_result_1;
  wire       [0:0]    Axi4Incr_sizeValue_1;
  wire       [11:0]   Axi4Incr_alignMask_1;
  wire       [11:0]   Axi4Incr_base_1;
  wire       [11:0]   Axi4Incr_baseIncr_1;
  reg        [1:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [1:0]    Axi4Incr_wrapCase_1;
  wire                when_Axi4_transmission_l174;
  wire                when_Axi4_transmission_l177;
  reg                 regLast;
  wire                when_Axi4_transmission_l182;
  wire                when_Axi4_transmission_l184;
  wire                when_Axi4_transmission_l189;
  wire                when_Axi4_transmission_l191;

  assign _zz_rFireCounter_valueNext_1 = rFireCounter_willIncrement;
  assign _zz_rFireCounter_valueNext = {12'd0, _zz_rFireCounter_valueNext_1};
  assign _zz_regAwAddr = axiSignal_aw_payload_addr;
  assign _zz__zz_1 = (regAwAddr + 12'h0);
  assign _zz__zz_regVec_0_1 = (regAwAddr + 12'h0);
  assign _zz_Axi4Incr_base_1 = regAwAddr[11 : 0];
  assign _zz_Axi4Incr_base = _zz_Axi4Incr_base_1;
  assign _zz_Axi4Incr_baseIncr = {11'd0, Axi4Incr_sizeValue};
  assign _zz_regArAddr = axiSignal_ar_payload_addr;
  assign _zz_axiSignal_r_payload_data_1 = (regArAddr + 12'h0);
  assign _zz_Axi4Incr_base_1_2 = regArAddr[11 : 0];
  assign _zz_Axi4Incr_base_1_1 = _zz_Axi4Incr_base_1_2;
  assign _zz_Axi4Incr_baseIncr_1 = {11'd0, Axi4Incr_sizeValue_1};
  assign _zz_when_Axi4_transmission_l177 = {5'd0, regArLen};
  assign _zz_when_Axi4_transmission_l182_1 = (regArLen - 8'h01);
  assign _zz_when_Axi4_transmission_l182 = {5'd0, _zz_when_Axi4_transmission_l182_1};
  always @(*) begin
    case(_zz__zz_regVec_0_1)
      12'b000000000000 : begin
        _zz__zz_regVec_0 = regVec_0;
      end
      12'b000000000001 : begin
        _zz__zz_regVec_0 = regVec_1;
      end
      12'b000000000010 : begin
        _zz__zz_regVec_0 = regVec_2;
      end
      12'b000000000011 : begin
        _zz__zz_regVec_0 = regVec_3;
      end
      12'b000000000100 : begin
        _zz__zz_regVec_0 = regVec_4;
      end
      12'b000000000101 : begin
        _zz__zz_regVec_0 = regVec_5;
      end
      12'b000000000110 : begin
        _zz__zz_regVec_0 = regVec_6;
      end
      12'b000000000111 : begin
        _zz__zz_regVec_0 = regVec_7;
      end
      12'b000000001000 : begin
        _zz__zz_regVec_0 = regVec_8;
      end
      12'b000000001001 : begin
        _zz__zz_regVec_0 = regVec_9;
      end
      12'b000000001010 : begin
        _zz__zz_regVec_0 = regVec_10;
      end
      12'b000000001011 : begin
        _zz__zz_regVec_0 = regVec_11;
      end
      12'b000000001100 : begin
        _zz__zz_regVec_0 = regVec_12;
      end
      12'b000000001101 : begin
        _zz__zz_regVec_0 = regVec_13;
      end
      12'b000000001110 : begin
        _zz__zz_regVec_0 = regVec_14;
      end
      12'b000000001111 : begin
        _zz__zz_regVec_0 = regVec_15;
      end
      12'b000000010000 : begin
        _zz__zz_regVec_0 = regVec_16;
      end
      12'b000000010001 : begin
        _zz__zz_regVec_0 = regVec_17;
      end
      12'b000000010010 : begin
        _zz__zz_regVec_0 = regVec_18;
      end
      12'b000000010011 : begin
        _zz__zz_regVec_0 = regVec_19;
      end
      12'b000000010100 : begin
        _zz__zz_regVec_0 = regVec_20;
      end
      12'b000000010101 : begin
        _zz__zz_regVec_0 = regVec_21;
      end
      12'b000000010110 : begin
        _zz__zz_regVec_0 = regVec_22;
      end
      12'b000000010111 : begin
        _zz__zz_regVec_0 = regVec_23;
      end
      12'b000000011000 : begin
        _zz__zz_regVec_0 = regVec_24;
      end
      12'b000000011001 : begin
        _zz__zz_regVec_0 = regVec_25;
      end
      12'b000000011010 : begin
        _zz__zz_regVec_0 = regVec_26;
      end
      12'b000000011011 : begin
        _zz__zz_regVec_0 = regVec_27;
      end
      12'b000000011100 : begin
        _zz__zz_regVec_0 = regVec_28;
      end
      12'b000000011101 : begin
        _zz__zz_regVec_0 = regVec_29;
      end
      12'b000000011110 : begin
        _zz__zz_regVec_0 = regVec_30;
      end
      12'b000000011111 : begin
        _zz__zz_regVec_0 = regVec_31;
      end
      12'b000000100000 : begin
        _zz__zz_regVec_0 = regVec_32;
      end
      12'b000000100001 : begin
        _zz__zz_regVec_0 = regVec_33;
      end
      12'b000000100010 : begin
        _zz__zz_regVec_0 = regVec_34;
      end
      12'b000000100011 : begin
        _zz__zz_regVec_0 = regVec_35;
      end
      12'b000000100100 : begin
        _zz__zz_regVec_0 = regVec_36;
      end
      12'b000000100101 : begin
        _zz__zz_regVec_0 = regVec_37;
      end
      12'b000000100110 : begin
        _zz__zz_regVec_0 = regVec_38;
      end
      12'b000000100111 : begin
        _zz__zz_regVec_0 = regVec_39;
      end
      12'b000000101000 : begin
        _zz__zz_regVec_0 = regVec_40;
      end
      12'b000000101001 : begin
        _zz__zz_regVec_0 = regVec_41;
      end
      12'b000000101010 : begin
        _zz__zz_regVec_0 = regVec_42;
      end
      12'b000000101011 : begin
        _zz__zz_regVec_0 = regVec_43;
      end
      12'b000000101100 : begin
        _zz__zz_regVec_0 = regVec_44;
      end
      12'b000000101101 : begin
        _zz__zz_regVec_0 = regVec_45;
      end
      12'b000000101110 : begin
        _zz__zz_regVec_0 = regVec_46;
      end
      12'b000000101111 : begin
        _zz__zz_regVec_0 = regVec_47;
      end
      12'b000000110000 : begin
        _zz__zz_regVec_0 = regVec_48;
      end
      12'b000000110001 : begin
        _zz__zz_regVec_0 = regVec_49;
      end
      12'b000000110010 : begin
        _zz__zz_regVec_0 = regVec_50;
      end
      12'b000000110011 : begin
        _zz__zz_regVec_0 = regVec_51;
      end
      12'b000000110100 : begin
        _zz__zz_regVec_0 = regVec_52;
      end
      12'b000000110101 : begin
        _zz__zz_regVec_0 = regVec_53;
      end
      12'b000000110110 : begin
        _zz__zz_regVec_0 = regVec_54;
      end
      12'b000000110111 : begin
        _zz__zz_regVec_0 = regVec_55;
      end
      12'b000000111000 : begin
        _zz__zz_regVec_0 = regVec_56;
      end
      12'b000000111001 : begin
        _zz__zz_regVec_0 = regVec_57;
      end
      12'b000000111010 : begin
        _zz__zz_regVec_0 = regVec_58;
      end
      12'b000000111011 : begin
        _zz__zz_regVec_0 = regVec_59;
      end
      12'b000000111100 : begin
        _zz__zz_regVec_0 = regVec_60;
      end
      12'b000000111101 : begin
        _zz__zz_regVec_0 = regVec_61;
      end
      12'b000000111110 : begin
        _zz__zz_regVec_0 = regVec_62;
      end
      12'b000000111111 : begin
        _zz__zz_regVec_0 = regVec_63;
      end
      12'b000001000000 : begin
        _zz__zz_regVec_0 = regVec_64;
      end
      12'b000001000001 : begin
        _zz__zz_regVec_0 = regVec_65;
      end
      12'b000001000010 : begin
        _zz__zz_regVec_0 = regVec_66;
      end
      12'b000001000011 : begin
        _zz__zz_regVec_0 = regVec_67;
      end
      12'b000001000100 : begin
        _zz__zz_regVec_0 = regVec_68;
      end
      12'b000001000101 : begin
        _zz__zz_regVec_0 = regVec_69;
      end
      12'b000001000110 : begin
        _zz__zz_regVec_0 = regVec_70;
      end
      12'b000001000111 : begin
        _zz__zz_regVec_0 = regVec_71;
      end
      12'b000001001000 : begin
        _zz__zz_regVec_0 = regVec_72;
      end
      12'b000001001001 : begin
        _zz__zz_regVec_0 = regVec_73;
      end
      12'b000001001010 : begin
        _zz__zz_regVec_0 = regVec_74;
      end
      12'b000001001011 : begin
        _zz__zz_regVec_0 = regVec_75;
      end
      12'b000001001100 : begin
        _zz__zz_regVec_0 = regVec_76;
      end
      12'b000001001101 : begin
        _zz__zz_regVec_0 = regVec_77;
      end
      12'b000001001110 : begin
        _zz__zz_regVec_0 = regVec_78;
      end
      12'b000001001111 : begin
        _zz__zz_regVec_0 = regVec_79;
      end
      12'b000001010000 : begin
        _zz__zz_regVec_0 = regVec_80;
      end
      12'b000001010001 : begin
        _zz__zz_regVec_0 = regVec_81;
      end
      12'b000001010010 : begin
        _zz__zz_regVec_0 = regVec_82;
      end
      12'b000001010011 : begin
        _zz__zz_regVec_0 = regVec_83;
      end
      12'b000001010100 : begin
        _zz__zz_regVec_0 = regVec_84;
      end
      12'b000001010101 : begin
        _zz__zz_regVec_0 = regVec_85;
      end
      12'b000001010110 : begin
        _zz__zz_regVec_0 = regVec_86;
      end
      12'b000001010111 : begin
        _zz__zz_regVec_0 = regVec_87;
      end
      12'b000001011000 : begin
        _zz__zz_regVec_0 = regVec_88;
      end
      12'b000001011001 : begin
        _zz__zz_regVec_0 = regVec_89;
      end
      12'b000001011010 : begin
        _zz__zz_regVec_0 = regVec_90;
      end
      12'b000001011011 : begin
        _zz__zz_regVec_0 = regVec_91;
      end
      12'b000001011100 : begin
        _zz__zz_regVec_0 = regVec_92;
      end
      12'b000001011101 : begin
        _zz__zz_regVec_0 = regVec_93;
      end
      12'b000001011110 : begin
        _zz__zz_regVec_0 = regVec_94;
      end
      12'b000001011111 : begin
        _zz__zz_regVec_0 = regVec_95;
      end
      12'b000001100000 : begin
        _zz__zz_regVec_0 = regVec_96;
      end
      12'b000001100001 : begin
        _zz__zz_regVec_0 = regVec_97;
      end
      12'b000001100010 : begin
        _zz__zz_regVec_0 = regVec_98;
      end
      12'b000001100011 : begin
        _zz__zz_regVec_0 = regVec_99;
      end
      12'b000001100100 : begin
        _zz__zz_regVec_0 = regVec_100;
      end
      12'b000001100101 : begin
        _zz__zz_regVec_0 = regVec_101;
      end
      12'b000001100110 : begin
        _zz__zz_regVec_0 = regVec_102;
      end
      12'b000001100111 : begin
        _zz__zz_regVec_0 = regVec_103;
      end
      12'b000001101000 : begin
        _zz__zz_regVec_0 = regVec_104;
      end
      12'b000001101001 : begin
        _zz__zz_regVec_0 = regVec_105;
      end
      12'b000001101010 : begin
        _zz__zz_regVec_0 = regVec_106;
      end
      12'b000001101011 : begin
        _zz__zz_regVec_0 = regVec_107;
      end
      12'b000001101100 : begin
        _zz__zz_regVec_0 = regVec_108;
      end
      12'b000001101101 : begin
        _zz__zz_regVec_0 = regVec_109;
      end
      12'b000001101110 : begin
        _zz__zz_regVec_0 = regVec_110;
      end
      12'b000001101111 : begin
        _zz__zz_regVec_0 = regVec_111;
      end
      12'b000001110000 : begin
        _zz__zz_regVec_0 = regVec_112;
      end
      12'b000001110001 : begin
        _zz__zz_regVec_0 = regVec_113;
      end
      12'b000001110010 : begin
        _zz__zz_regVec_0 = regVec_114;
      end
      12'b000001110011 : begin
        _zz__zz_regVec_0 = regVec_115;
      end
      12'b000001110100 : begin
        _zz__zz_regVec_0 = regVec_116;
      end
      12'b000001110101 : begin
        _zz__zz_regVec_0 = regVec_117;
      end
      12'b000001110110 : begin
        _zz__zz_regVec_0 = regVec_118;
      end
      12'b000001110111 : begin
        _zz__zz_regVec_0 = regVec_119;
      end
      12'b000001111000 : begin
        _zz__zz_regVec_0 = regVec_120;
      end
      12'b000001111001 : begin
        _zz__zz_regVec_0 = regVec_121;
      end
      12'b000001111010 : begin
        _zz__zz_regVec_0 = regVec_122;
      end
      12'b000001111011 : begin
        _zz__zz_regVec_0 = regVec_123;
      end
      12'b000001111100 : begin
        _zz__zz_regVec_0 = regVec_124;
      end
      12'b000001111101 : begin
        _zz__zz_regVec_0 = regVec_125;
      end
      12'b000001111110 : begin
        _zz__zz_regVec_0 = regVec_126;
      end
      12'b000001111111 : begin
        _zz__zz_regVec_0 = regVec_127;
      end
      12'b000010000000 : begin
        _zz__zz_regVec_0 = regVec_128;
      end
      12'b000010000001 : begin
        _zz__zz_regVec_0 = regVec_129;
      end
      12'b000010000010 : begin
        _zz__zz_regVec_0 = regVec_130;
      end
      12'b000010000011 : begin
        _zz__zz_regVec_0 = regVec_131;
      end
      12'b000010000100 : begin
        _zz__zz_regVec_0 = regVec_132;
      end
      12'b000010000101 : begin
        _zz__zz_regVec_0 = regVec_133;
      end
      12'b000010000110 : begin
        _zz__zz_regVec_0 = regVec_134;
      end
      12'b000010000111 : begin
        _zz__zz_regVec_0 = regVec_135;
      end
      12'b000010001000 : begin
        _zz__zz_regVec_0 = regVec_136;
      end
      12'b000010001001 : begin
        _zz__zz_regVec_0 = regVec_137;
      end
      12'b000010001010 : begin
        _zz__zz_regVec_0 = regVec_138;
      end
      12'b000010001011 : begin
        _zz__zz_regVec_0 = regVec_139;
      end
      12'b000010001100 : begin
        _zz__zz_regVec_0 = regVec_140;
      end
      12'b000010001101 : begin
        _zz__zz_regVec_0 = regVec_141;
      end
      12'b000010001110 : begin
        _zz__zz_regVec_0 = regVec_142;
      end
      12'b000010001111 : begin
        _zz__zz_regVec_0 = regVec_143;
      end
      12'b000010010000 : begin
        _zz__zz_regVec_0 = regVec_144;
      end
      12'b000010010001 : begin
        _zz__zz_regVec_0 = regVec_145;
      end
      12'b000010010010 : begin
        _zz__zz_regVec_0 = regVec_146;
      end
      12'b000010010011 : begin
        _zz__zz_regVec_0 = regVec_147;
      end
      12'b000010010100 : begin
        _zz__zz_regVec_0 = regVec_148;
      end
      12'b000010010101 : begin
        _zz__zz_regVec_0 = regVec_149;
      end
      12'b000010010110 : begin
        _zz__zz_regVec_0 = regVec_150;
      end
      12'b000010010111 : begin
        _zz__zz_regVec_0 = regVec_151;
      end
      12'b000010011000 : begin
        _zz__zz_regVec_0 = regVec_152;
      end
      12'b000010011001 : begin
        _zz__zz_regVec_0 = regVec_153;
      end
      12'b000010011010 : begin
        _zz__zz_regVec_0 = regVec_154;
      end
      12'b000010011011 : begin
        _zz__zz_regVec_0 = regVec_155;
      end
      12'b000010011100 : begin
        _zz__zz_regVec_0 = regVec_156;
      end
      12'b000010011101 : begin
        _zz__zz_regVec_0 = regVec_157;
      end
      12'b000010011110 : begin
        _zz__zz_regVec_0 = regVec_158;
      end
      12'b000010011111 : begin
        _zz__zz_regVec_0 = regVec_159;
      end
      12'b000010100000 : begin
        _zz__zz_regVec_0 = regVec_160;
      end
      12'b000010100001 : begin
        _zz__zz_regVec_0 = regVec_161;
      end
      12'b000010100010 : begin
        _zz__zz_regVec_0 = regVec_162;
      end
      12'b000010100011 : begin
        _zz__zz_regVec_0 = regVec_163;
      end
      12'b000010100100 : begin
        _zz__zz_regVec_0 = regVec_164;
      end
      12'b000010100101 : begin
        _zz__zz_regVec_0 = regVec_165;
      end
      12'b000010100110 : begin
        _zz__zz_regVec_0 = regVec_166;
      end
      12'b000010100111 : begin
        _zz__zz_regVec_0 = regVec_167;
      end
      12'b000010101000 : begin
        _zz__zz_regVec_0 = regVec_168;
      end
      12'b000010101001 : begin
        _zz__zz_regVec_0 = regVec_169;
      end
      12'b000010101010 : begin
        _zz__zz_regVec_0 = regVec_170;
      end
      12'b000010101011 : begin
        _zz__zz_regVec_0 = regVec_171;
      end
      12'b000010101100 : begin
        _zz__zz_regVec_0 = regVec_172;
      end
      12'b000010101101 : begin
        _zz__zz_regVec_0 = regVec_173;
      end
      12'b000010101110 : begin
        _zz__zz_regVec_0 = regVec_174;
      end
      12'b000010101111 : begin
        _zz__zz_regVec_0 = regVec_175;
      end
      12'b000010110000 : begin
        _zz__zz_regVec_0 = regVec_176;
      end
      12'b000010110001 : begin
        _zz__zz_regVec_0 = regVec_177;
      end
      12'b000010110010 : begin
        _zz__zz_regVec_0 = regVec_178;
      end
      12'b000010110011 : begin
        _zz__zz_regVec_0 = regVec_179;
      end
      12'b000010110100 : begin
        _zz__zz_regVec_0 = regVec_180;
      end
      12'b000010110101 : begin
        _zz__zz_regVec_0 = regVec_181;
      end
      12'b000010110110 : begin
        _zz__zz_regVec_0 = regVec_182;
      end
      12'b000010110111 : begin
        _zz__zz_regVec_0 = regVec_183;
      end
      12'b000010111000 : begin
        _zz__zz_regVec_0 = regVec_184;
      end
      12'b000010111001 : begin
        _zz__zz_regVec_0 = regVec_185;
      end
      12'b000010111010 : begin
        _zz__zz_regVec_0 = regVec_186;
      end
      12'b000010111011 : begin
        _zz__zz_regVec_0 = regVec_187;
      end
      12'b000010111100 : begin
        _zz__zz_regVec_0 = regVec_188;
      end
      12'b000010111101 : begin
        _zz__zz_regVec_0 = regVec_189;
      end
      12'b000010111110 : begin
        _zz__zz_regVec_0 = regVec_190;
      end
      12'b000010111111 : begin
        _zz__zz_regVec_0 = regVec_191;
      end
      12'b000011000000 : begin
        _zz__zz_regVec_0 = regVec_192;
      end
      12'b000011000001 : begin
        _zz__zz_regVec_0 = regVec_193;
      end
      12'b000011000010 : begin
        _zz__zz_regVec_0 = regVec_194;
      end
      12'b000011000011 : begin
        _zz__zz_regVec_0 = regVec_195;
      end
      12'b000011000100 : begin
        _zz__zz_regVec_0 = regVec_196;
      end
      12'b000011000101 : begin
        _zz__zz_regVec_0 = regVec_197;
      end
      12'b000011000110 : begin
        _zz__zz_regVec_0 = regVec_198;
      end
      12'b000011000111 : begin
        _zz__zz_regVec_0 = regVec_199;
      end
      12'b000011001000 : begin
        _zz__zz_regVec_0 = regVec_200;
      end
      12'b000011001001 : begin
        _zz__zz_regVec_0 = regVec_201;
      end
      12'b000011001010 : begin
        _zz__zz_regVec_0 = regVec_202;
      end
      12'b000011001011 : begin
        _zz__zz_regVec_0 = regVec_203;
      end
      12'b000011001100 : begin
        _zz__zz_regVec_0 = regVec_204;
      end
      12'b000011001101 : begin
        _zz__zz_regVec_0 = regVec_205;
      end
      12'b000011001110 : begin
        _zz__zz_regVec_0 = regVec_206;
      end
      12'b000011001111 : begin
        _zz__zz_regVec_0 = regVec_207;
      end
      12'b000011010000 : begin
        _zz__zz_regVec_0 = regVec_208;
      end
      12'b000011010001 : begin
        _zz__zz_regVec_0 = regVec_209;
      end
      12'b000011010010 : begin
        _zz__zz_regVec_0 = regVec_210;
      end
      12'b000011010011 : begin
        _zz__zz_regVec_0 = regVec_211;
      end
      12'b000011010100 : begin
        _zz__zz_regVec_0 = regVec_212;
      end
      12'b000011010101 : begin
        _zz__zz_regVec_0 = regVec_213;
      end
      12'b000011010110 : begin
        _zz__zz_regVec_0 = regVec_214;
      end
      12'b000011010111 : begin
        _zz__zz_regVec_0 = regVec_215;
      end
      12'b000011011000 : begin
        _zz__zz_regVec_0 = regVec_216;
      end
      12'b000011011001 : begin
        _zz__zz_regVec_0 = regVec_217;
      end
      12'b000011011010 : begin
        _zz__zz_regVec_0 = regVec_218;
      end
      12'b000011011011 : begin
        _zz__zz_regVec_0 = regVec_219;
      end
      12'b000011011100 : begin
        _zz__zz_regVec_0 = regVec_220;
      end
      12'b000011011101 : begin
        _zz__zz_regVec_0 = regVec_221;
      end
      12'b000011011110 : begin
        _zz__zz_regVec_0 = regVec_222;
      end
      12'b000011011111 : begin
        _zz__zz_regVec_0 = regVec_223;
      end
      12'b000011100000 : begin
        _zz__zz_regVec_0 = regVec_224;
      end
      12'b000011100001 : begin
        _zz__zz_regVec_0 = regVec_225;
      end
      12'b000011100010 : begin
        _zz__zz_regVec_0 = regVec_226;
      end
      12'b000011100011 : begin
        _zz__zz_regVec_0 = regVec_227;
      end
      12'b000011100100 : begin
        _zz__zz_regVec_0 = regVec_228;
      end
      12'b000011100101 : begin
        _zz__zz_regVec_0 = regVec_229;
      end
      12'b000011100110 : begin
        _zz__zz_regVec_0 = regVec_230;
      end
      12'b000011100111 : begin
        _zz__zz_regVec_0 = regVec_231;
      end
      12'b000011101000 : begin
        _zz__zz_regVec_0 = regVec_232;
      end
      12'b000011101001 : begin
        _zz__zz_regVec_0 = regVec_233;
      end
      12'b000011101010 : begin
        _zz__zz_regVec_0 = regVec_234;
      end
      12'b000011101011 : begin
        _zz__zz_regVec_0 = regVec_235;
      end
      12'b000011101100 : begin
        _zz__zz_regVec_0 = regVec_236;
      end
      12'b000011101101 : begin
        _zz__zz_regVec_0 = regVec_237;
      end
      12'b000011101110 : begin
        _zz__zz_regVec_0 = regVec_238;
      end
      12'b000011101111 : begin
        _zz__zz_regVec_0 = regVec_239;
      end
      12'b000011110000 : begin
        _zz__zz_regVec_0 = regVec_240;
      end
      12'b000011110001 : begin
        _zz__zz_regVec_0 = regVec_241;
      end
      12'b000011110010 : begin
        _zz__zz_regVec_0 = regVec_242;
      end
      12'b000011110011 : begin
        _zz__zz_regVec_0 = regVec_243;
      end
      12'b000011110100 : begin
        _zz__zz_regVec_0 = regVec_244;
      end
      12'b000011110101 : begin
        _zz__zz_regVec_0 = regVec_245;
      end
      12'b000011110110 : begin
        _zz__zz_regVec_0 = regVec_246;
      end
      12'b000011110111 : begin
        _zz__zz_regVec_0 = regVec_247;
      end
      12'b000011111000 : begin
        _zz__zz_regVec_0 = regVec_248;
      end
      12'b000011111001 : begin
        _zz__zz_regVec_0 = regVec_249;
      end
      12'b000011111010 : begin
        _zz__zz_regVec_0 = regVec_250;
      end
      12'b000011111011 : begin
        _zz__zz_regVec_0 = regVec_251;
      end
      12'b000011111100 : begin
        _zz__zz_regVec_0 = regVec_252;
      end
      12'b000011111101 : begin
        _zz__zz_regVec_0 = regVec_253;
      end
      12'b000011111110 : begin
        _zz__zz_regVec_0 = regVec_254;
      end
      12'b000011111111 : begin
        _zz__zz_regVec_0 = regVec_255;
      end
      12'b000100000000 : begin
        _zz__zz_regVec_0 = regVec_256;
      end
      12'b000100000001 : begin
        _zz__zz_regVec_0 = regVec_257;
      end
      12'b000100000010 : begin
        _zz__zz_regVec_0 = regVec_258;
      end
      12'b000100000011 : begin
        _zz__zz_regVec_0 = regVec_259;
      end
      12'b000100000100 : begin
        _zz__zz_regVec_0 = regVec_260;
      end
      12'b000100000101 : begin
        _zz__zz_regVec_0 = regVec_261;
      end
      12'b000100000110 : begin
        _zz__zz_regVec_0 = regVec_262;
      end
      12'b000100000111 : begin
        _zz__zz_regVec_0 = regVec_263;
      end
      12'b000100001000 : begin
        _zz__zz_regVec_0 = regVec_264;
      end
      12'b000100001001 : begin
        _zz__zz_regVec_0 = regVec_265;
      end
      12'b000100001010 : begin
        _zz__zz_regVec_0 = regVec_266;
      end
      12'b000100001011 : begin
        _zz__zz_regVec_0 = regVec_267;
      end
      12'b000100001100 : begin
        _zz__zz_regVec_0 = regVec_268;
      end
      12'b000100001101 : begin
        _zz__zz_regVec_0 = regVec_269;
      end
      12'b000100001110 : begin
        _zz__zz_regVec_0 = regVec_270;
      end
      12'b000100001111 : begin
        _zz__zz_regVec_0 = regVec_271;
      end
      12'b000100010000 : begin
        _zz__zz_regVec_0 = regVec_272;
      end
      12'b000100010001 : begin
        _zz__zz_regVec_0 = regVec_273;
      end
      12'b000100010010 : begin
        _zz__zz_regVec_0 = regVec_274;
      end
      12'b000100010011 : begin
        _zz__zz_regVec_0 = regVec_275;
      end
      12'b000100010100 : begin
        _zz__zz_regVec_0 = regVec_276;
      end
      12'b000100010101 : begin
        _zz__zz_regVec_0 = regVec_277;
      end
      12'b000100010110 : begin
        _zz__zz_regVec_0 = regVec_278;
      end
      12'b000100010111 : begin
        _zz__zz_regVec_0 = regVec_279;
      end
      12'b000100011000 : begin
        _zz__zz_regVec_0 = regVec_280;
      end
      12'b000100011001 : begin
        _zz__zz_regVec_0 = regVec_281;
      end
      12'b000100011010 : begin
        _zz__zz_regVec_0 = regVec_282;
      end
      12'b000100011011 : begin
        _zz__zz_regVec_0 = regVec_283;
      end
      12'b000100011100 : begin
        _zz__zz_regVec_0 = regVec_284;
      end
      12'b000100011101 : begin
        _zz__zz_regVec_0 = regVec_285;
      end
      12'b000100011110 : begin
        _zz__zz_regVec_0 = regVec_286;
      end
      12'b000100011111 : begin
        _zz__zz_regVec_0 = regVec_287;
      end
      12'b000100100000 : begin
        _zz__zz_regVec_0 = regVec_288;
      end
      12'b000100100001 : begin
        _zz__zz_regVec_0 = regVec_289;
      end
      12'b000100100010 : begin
        _zz__zz_regVec_0 = regVec_290;
      end
      12'b000100100011 : begin
        _zz__zz_regVec_0 = regVec_291;
      end
      12'b000100100100 : begin
        _zz__zz_regVec_0 = regVec_292;
      end
      12'b000100100101 : begin
        _zz__zz_regVec_0 = regVec_293;
      end
      12'b000100100110 : begin
        _zz__zz_regVec_0 = regVec_294;
      end
      12'b000100100111 : begin
        _zz__zz_regVec_0 = regVec_295;
      end
      12'b000100101000 : begin
        _zz__zz_regVec_0 = regVec_296;
      end
      12'b000100101001 : begin
        _zz__zz_regVec_0 = regVec_297;
      end
      12'b000100101010 : begin
        _zz__zz_regVec_0 = regVec_298;
      end
      12'b000100101011 : begin
        _zz__zz_regVec_0 = regVec_299;
      end
      12'b000100101100 : begin
        _zz__zz_regVec_0 = regVec_300;
      end
      12'b000100101101 : begin
        _zz__zz_regVec_0 = regVec_301;
      end
      12'b000100101110 : begin
        _zz__zz_regVec_0 = regVec_302;
      end
      12'b000100101111 : begin
        _zz__zz_regVec_0 = regVec_303;
      end
      12'b000100110000 : begin
        _zz__zz_regVec_0 = regVec_304;
      end
      12'b000100110001 : begin
        _zz__zz_regVec_0 = regVec_305;
      end
      12'b000100110010 : begin
        _zz__zz_regVec_0 = regVec_306;
      end
      12'b000100110011 : begin
        _zz__zz_regVec_0 = regVec_307;
      end
      12'b000100110100 : begin
        _zz__zz_regVec_0 = regVec_308;
      end
      12'b000100110101 : begin
        _zz__zz_regVec_0 = regVec_309;
      end
      12'b000100110110 : begin
        _zz__zz_regVec_0 = regVec_310;
      end
      12'b000100110111 : begin
        _zz__zz_regVec_0 = regVec_311;
      end
      12'b000100111000 : begin
        _zz__zz_regVec_0 = regVec_312;
      end
      12'b000100111001 : begin
        _zz__zz_regVec_0 = regVec_313;
      end
      12'b000100111010 : begin
        _zz__zz_regVec_0 = regVec_314;
      end
      12'b000100111011 : begin
        _zz__zz_regVec_0 = regVec_315;
      end
      12'b000100111100 : begin
        _zz__zz_regVec_0 = regVec_316;
      end
      12'b000100111101 : begin
        _zz__zz_regVec_0 = regVec_317;
      end
      12'b000100111110 : begin
        _zz__zz_regVec_0 = regVec_318;
      end
      12'b000100111111 : begin
        _zz__zz_regVec_0 = regVec_319;
      end
      12'b000101000000 : begin
        _zz__zz_regVec_0 = regVec_320;
      end
      12'b000101000001 : begin
        _zz__zz_regVec_0 = regVec_321;
      end
      12'b000101000010 : begin
        _zz__zz_regVec_0 = regVec_322;
      end
      12'b000101000011 : begin
        _zz__zz_regVec_0 = regVec_323;
      end
      12'b000101000100 : begin
        _zz__zz_regVec_0 = regVec_324;
      end
      12'b000101000101 : begin
        _zz__zz_regVec_0 = regVec_325;
      end
      12'b000101000110 : begin
        _zz__zz_regVec_0 = regVec_326;
      end
      12'b000101000111 : begin
        _zz__zz_regVec_0 = regVec_327;
      end
      12'b000101001000 : begin
        _zz__zz_regVec_0 = regVec_328;
      end
      12'b000101001001 : begin
        _zz__zz_regVec_0 = regVec_329;
      end
      12'b000101001010 : begin
        _zz__zz_regVec_0 = regVec_330;
      end
      12'b000101001011 : begin
        _zz__zz_regVec_0 = regVec_331;
      end
      12'b000101001100 : begin
        _zz__zz_regVec_0 = regVec_332;
      end
      12'b000101001101 : begin
        _zz__zz_regVec_0 = regVec_333;
      end
      12'b000101001110 : begin
        _zz__zz_regVec_0 = regVec_334;
      end
      12'b000101001111 : begin
        _zz__zz_regVec_0 = regVec_335;
      end
      12'b000101010000 : begin
        _zz__zz_regVec_0 = regVec_336;
      end
      12'b000101010001 : begin
        _zz__zz_regVec_0 = regVec_337;
      end
      12'b000101010010 : begin
        _zz__zz_regVec_0 = regVec_338;
      end
      12'b000101010011 : begin
        _zz__zz_regVec_0 = regVec_339;
      end
      12'b000101010100 : begin
        _zz__zz_regVec_0 = regVec_340;
      end
      12'b000101010101 : begin
        _zz__zz_regVec_0 = regVec_341;
      end
      12'b000101010110 : begin
        _zz__zz_regVec_0 = regVec_342;
      end
      12'b000101010111 : begin
        _zz__zz_regVec_0 = regVec_343;
      end
      12'b000101011000 : begin
        _zz__zz_regVec_0 = regVec_344;
      end
      12'b000101011001 : begin
        _zz__zz_regVec_0 = regVec_345;
      end
      12'b000101011010 : begin
        _zz__zz_regVec_0 = regVec_346;
      end
      12'b000101011011 : begin
        _zz__zz_regVec_0 = regVec_347;
      end
      12'b000101011100 : begin
        _zz__zz_regVec_0 = regVec_348;
      end
      12'b000101011101 : begin
        _zz__zz_regVec_0 = regVec_349;
      end
      12'b000101011110 : begin
        _zz__zz_regVec_0 = regVec_350;
      end
      12'b000101011111 : begin
        _zz__zz_regVec_0 = regVec_351;
      end
      12'b000101100000 : begin
        _zz__zz_regVec_0 = regVec_352;
      end
      12'b000101100001 : begin
        _zz__zz_regVec_0 = regVec_353;
      end
      12'b000101100010 : begin
        _zz__zz_regVec_0 = regVec_354;
      end
      12'b000101100011 : begin
        _zz__zz_regVec_0 = regVec_355;
      end
      12'b000101100100 : begin
        _zz__zz_regVec_0 = regVec_356;
      end
      12'b000101100101 : begin
        _zz__zz_regVec_0 = regVec_357;
      end
      12'b000101100110 : begin
        _zz__zz_regVec_0 = regVec_358;
      end
      12'b000101100111 : begin
        _zz__zz_regVec_0 = regVec_359;
      end
      12'b000101101000 : begin
        _zz__zz_regVec_0 = regVec_360;
      end
      12'b000101101001 : begin
        _zz__zz_regVec_0 = regVec_361;
      end
      12'b000101101010 : begin
        _zz__zz_regVec_0 = regVec_362;
      end
      12'b000101101011 : begin
        _zz__zz_regVec_0 = regVec_363;
      end
      12'b000101101100 : begin
        _zz__zz_regVec_0 = regVec_364;
      end
      12'b000101101101 : begin
        _zz__zz_regVec_0 = regVec_365;
      end
      12'b000101101110 : begin
        _zz__zz_regVec_0 = regVec_366;
      end
      12'b000101101111 : begin
        _zz__zz_regVec_0 = regVec_367;
      end
      12'b000101110000 : begin
        _zz__zz_regVec_0 = regVec_368;
      end
      12'b000101110001 : begin
        _zz__zz_regVec_0 = regVec_369;
      end
      12'b000101110010 : begin
        _zz__zz_regVec_0 = regVec_370;
      end
      12'b000101110011 : begin
        _zz__zz_regVec_0 = regVec_371;
      end
      12'b000101110100 : begin
        _zz__zz_regVec_0 = regVec_372;
      end
      12'b000101110101 : begin
        _zz__zz_regVec_0 = regVec_373;
      end
      12'b000101110110 : begin
        _zz__zz_regVec_0 = regVec_374;
      end
      12'b000101110111 : begin
        _zz__zz_regVec_0 = regVec_375;
      end
      12'b000101111000 : begin
        _zz__zz_regVec_0 = regVec_376;
      end
      12'b000101111001 : begin
        _zz__zz_regVec_0 = regVec_377;
      end
      12'b000101111010 : begin
        _zz__zz_regVec_0 = regVec_378;
      end
      12'b000101111011 : begin
        _zz__zz_regVec_0 = regVec_379;
      end
      12'b000101111100 : begin
        _zz__zz_regVec_0 = regVec_380;
      end
      12'b000101111101 : begin
        _zz__zz_regVec_0 = regVec_381;
      end
      12'b000101111110 : begin
        _zz__zz_regVec_0 = regVec_382;
      end
      12'b000101111111 : begin
        _zz__zz_regVec_0 = regVec_383;
      end
      12'b000110000000 : begin
        _zz__zz_regVec_0 = regVec_384;
      end
      12'b000110000001 : begin
        _zz__zz_regVec_0 = regVec_385;
      end
      12'b000110000010 : begin
        _zz__zz_regVec_0 = regVec_386;
      end
      12'b000110000011 : begin
        _zz__zz_regVec_0 = regVec_387;
      end
      12'b000110000100 : begin
        _zz__zz_regVec_0 = regVec_388;
      end
      12'b000110000101 : begin
        _zz__zz_regVec_0 = regVec_389;
      end
      12'b000110000110 : begin
        _zz__zz_regVec_0 = regVec_390;
      end
      12'b000110000111 : begin
        _zz__zz_regVec_0 = regVec_391;
      end
      12'b000110001000 : begin
        _zz__zz_regVec_0 = regVec_392;
      end
      12'b000110001001 : begin
        _zz__zz_regVec_0 = regVec_393;
      end
      12'b000110001010 : begin
        _zz__zz_regVec_0 = regVec_394;
      end
      12'b000110001011 : begin
        _zz__zz_regVec_0 = regVec_395;
      end
      12'b000110001100 : begin
        _zz__zz_regVec_0 = regVec_396;
      end
      12'b000110001101 : begin
        _zz__zz_regVec_0 = regVec_397;
      end
      12'b000110001110 : begin
        _zz__zz_regVec_0 = regVec_398;
      end
      12'b000110001111 : begin
        _zz__zz_regVec_0 = regVec_399;
      end
      12'b000110010000 : begin
        _zz__zz_regVec_0 = regVec_400;
      end
      12'b000110010001 : begin
        _zz__zz_regVec_0 = regVec_401;
      end
      12'b000110010010 : begin
        _zz__zz_regVec_0 = regVec_402;
      end
      12'b000110010011 : begin
        _zz__zz_regVec_0 = regVec_403;
      end
      12'b000110010100 : begin
        _zz__zz_regVec_0 = regVec_404;
      end
      12'b000110010101 : begin
        _zz__zz_regVec_0 = regVec_405;
      end
      12'b000110010110 : begin
        _zz__zz_regVec_0 = regVec_406;
      end
      12'b000110010111 : begin
        _zz__zz_regVec_0 = regVec_407;
      end
      12'b000110011000 : begin
        _zz__zz_regVec_0 = regVec_408;
      end
      12'b000110011001 : begin
        _zz__zz_regVec_0 = regVec_409;
      end
      12'b000110011010 : begin
        _zz__zz_regVec_0 = regVec_410;
      end
      12'b000110011011 : begin
        _zz__zz_regVec_0 = regVec_411;
      end
      12'b000110011100 : begin
        _zz__zz_regVec_0 = regVec_412;
      end
      12'b000110011101 : begin
        _zz__zz_regVec_0 = regVec_413;
      end
      12'b000110011110 : begin
        _zz__zz_regVec_0 = regVec_414;
      end
      12'b000110011111 : begin
        _zz__zz_regVec_0 = regVec_415;
      end
      12'b000110100000 : begin
        _zz__zz_regVec_0 = regVec_416;
      end
      12'b000110100001 : begin
        _zz__zz_regVec_0 = regVec_417;
      end
      12'b000110100010 : begin
        _zz__zz_regVec_0 = regVec_418;
      end
      12'b000110100011 : begin
        _zz__zz_regVec_0 = regVec_419;
      end
      12'b000110100100 : begin
        _zz__zz_regVec_0 = regVec_420;
      end
      12'b000110100101 : begin
        _zz__zz_regVec_0 = regVec_421;
      end
      12'b000110100110 : begin
        _zz__zz_regVec_0 = regVec_422;
      end
      12'b000110100111 : begin
        _zz__zz_regVec_0 = regVec_423;
      end
      12'b000110101000 : begin
        _zz__zz_regVec_0 = regVec_424;
      end
      12'b000110101001 : begin
        _zz__zz_regVec_0 = regVec_425;
      end
      12'b000110101010 : begin
        _zz__zz_regVec_0 = regVec_426;
      end
      12'b000110101011 : begin
        _zz__zz_regVec_0 = regVec_427;
      end
      12'b000110101100 : begin
        _zz__zz_regVec_0 = regVec_428;
      end
      12'b000110101101 : begin
        _zz__zz_regVec_0 = regVec_429;
      end
      12'b000110101110 : begin
        _zz__zz_regVec_0 = regVec_430;
      end
      12'b000110101111 : begin
        _zz__zz_regVec_0 = regVec_431;
      end
      12'b000110110000 : begin
        _zz__zz_regVec_0 = regVec_432;
      end
      12'b000110110001 : begin
        _zz__zz_regVec_0 = regVec_433;
      end
      12'b000110110010 : begin
        _zz__zz_regVec_0 = regVec_434;
      end
      12'b000110110011 : begin
        _zz__zz_regVec_0 = regVec_435;
      end
      12'b000110110100 : begin
        _zz__zz_regVec_0 = regVec_436;
      end
      12'b000110110101 : begin
        _zz__zz_regVec_0 = regVec_437;
      end
      12'b000110110110 : begin
        _zz__zz_regVec_0 = regVec_438;
      end
      12'b000110110111 : begin
        _zz__zz_regVec_0 = regVec_439;
      end
      12'b000110111000 : begin
        _zz__zz_regVec_0 = regVec_440;
      end
      12'b000110111001 : begin
        _zz__zz_regVec_0 = regVec_441;
      end
      12'b000110111010 : begin
        _zz__zz_regVec_0 = regVec_442;
      end
      12'b000110111011 : begin
        _zz__zz_regVec_0 = regVec_443;
      end
      12'b000110111100 : begin
        _zz__zz_regVec_0 = regVec_444;
      end
      12'b000110111101 : begin
        _zz__zz_regVec_0 = regVec_445;
      end
      12'b000110111110 : begin
        _zz__zz_regVec_0 = regVec_446;
      end
      12'b000110111111 : begin
        _zz__zz_regVec_0 = regVec_447;
      end
      12'b000111000000 : begin
        _zz__zz_regVec_0 = regVec_448;
      end
      12'b000111000001 : begin
        _zz__zz_regVec_0 = regVec_449;
      end
      12'b000111000010 : begin
        _zz__zz_regVec_0 = regVec_450;
      end
      12'b000111000011 : begin
        _zz__zz_regVec_0 = regVec_451;
      end
      12'b000111000100 : begin
        _zz__zz_regVec_0 = regVec_452;
      end
      12'b000111000101 : begin
        _zz__zz_regVec_0 = regVec_453;
      end
      12'b000111000110 : begin
        _zz__zz_regVec_0 = regVec_454;
      end
      12'b000111000111 : begin
        _zz__zz_regVec_0 = regVec_455;
      end
      12'b000111001000 : begin
        _zz__zz_regVec_0 = regVec_456;
      end
      12'b000111001001 : begin
        _zz__zz_regVec_0 = regVec_457;
      end
      12'b000111001010 : begin
        _zz__zz_regVec_0 = regVec_458;
      end
      12'b000111001011 : begin
        _zz__zz_regVec_0 = regVec_459;
      end
      12'b000111001100 : begin
        _zz__zz_regVec_0 = regVec_460;
      end
      12'b000111001101 : begin
        _zz__zz_regVec_0 = regVec_461;
      end
      12'b000111001110 : begin
        _zz__zz_regVec_0 = regVec_462;
      end
      12'b000111001111 : begin
        _zz__zz_regVec_0 = regVec_463;
      end
      12'b000111010000 : begin
        _zz__zz_regVec_0 = regVec_464;
      end
      12'b000111010001 : begin
        _zz__zz_regVec_0 = regVec_465;
      end
      12'b000111010010 : begin
        _zz__zz_regVec_0 = regVec_466;
      end
      12'b000111010011 : begin
        _zz__zz_regVec_0 = regVec_467;
      end
      12'b000111010100 : begin
        _zz__zz_regVec_0 = regVec_468;
      end
      12'b000111010101 : begin
        _zz__zz_regVec_0 = regVec_469;
      end
      12'b000111010110 : begin
        _zz__zz_regVec_0 = regVec_470;
      end
      12'b000111010111 : begin
        _zz__zz_regVec_0 = regVec_471;
      end
      12'b000111011000 : begin
        _zz__zz_regVec_0 = regVec_472;
      end
      12'b000111011001 : begin
        _zz__zz_regVec_0 = regVec_473;
      end
      12'b000111011010 : begin
        _zz__zz_regVec_0 = regVec_474;
      end
      12'b000111011011 : begin
        _zz__zz_regVec_0 = regVec_475;
      end
      12'b000111011100 : begin
        _zz__zz_regVec_0 = regVec_476;
      end
      12'b000111011101 : begin
        _zz__zz_regVec_0 = regVec_477;
      end
      12'b000111011110 : begin
        _zz__zz_regVec_0 = regVec_478;
      end
      12'b000111011111 : begin
        _zz__zz_regVec_0 = regVec_479;
      end
      12'b000111100000 : begin
        _zz__zz_regVec_0 = regVec_480;
      end
      12'b000111100001 : begin
        _zz__zz_regVec_0 = regVec_481;
      end
      12'b000111100010 : begin
        _zz__zz_regVec_0 = regVec_482;
      end
      12'b000111100011 : begin
        _zz__zz_regVec_0 = regVec_483;
      end
      12'b000111100100 : begin
        _zz__zz_regVec_0 = regVec_484;
      end
      12'b000111100101 : begin
        _zz__zz_regVec_0 = regVec_485;
      end
      12'b000111100110 : begin
        _zz__zz_regVec_0 = regVec_486;
      end
      12'b000111100111 : begin
        _zz__zz_regVec_0 = regVec_487;
      end
      12'b000111101000 : begin
        _zz__zz_regVec_0 = regVec_488;
      end
      12'b000111101001 : begin
        _zz__zz_regVec_0 = regVec_489;
      end
      12'b000111101010 : begin
        _zz__zz_regVec_0 = regVec_490;
      end
      12'b000111101011 : begin
        _zz__zz_regVec_0 = regVec_491;
      end
      12'b000111101100 : begin
        _zz__zz_regVec_0 = regVec_492;
      end
      12'b000111101101 : begin
        _zz__zz_regVec_0 = regVec_493;
      end
      12'b000111101110 : begin
        _zz__zz_regVec_0 = regVec_494;
      end
      12'b000111101111 : begin
        _zz__zz_regVec_0 = regVec_495;
      end
      12'b000111110000 : begin
        _zz__zz_regVec_0 = regVec_496;
      end
      12'b000111110001 : begin
        _zz__zz_regVec_0 = regVec_497;
      end
      12'b000111110010 : begin
        _zz__zz_regVec_0 = regVec_498;
      end
      12'b000111110011 : begin
        _zz__zz_regVec_0 = regVec_499;
      end
      12'b000111110100 : begin
        _zz__zz_regVec_0 = regVec_500;
      end
      12'b000111110101 : begin
        _zz__zz_regVec_0 = regVec_501;
      end
      12'b000111110110 : begin
        _zz__zz_regVec_0 = regVec_502;
      end
      12'b000111110111 : begin
        _zz__zz_regVec_0 = regVec_503;
      end
      12'b000111111000 : begin
        _zz__zz_regVec_0 = regVec_504;
      end
      12'b000111111001 : begin
        _zz__zz_regVec_0 = regVec_505;
      end
      12'b000111111010 : begin
        _zz__zz_regVec_0 = regVec_506;
      end
      12'b000111111011 : begin
        _zz__zz_regVec_0 = regVec_507;
      end
      12'b000111111100 : begin
        _zz__zz_regVec_0 = regVec_508;
      end
      12'b000111111101 : begin
        _zz__zz_regVec_0 = regVec_509;
      end
      12'b000111111110 : begin
        _zz__zz_regVec_0 = regVec_510;
      end
      12'b000111111111 : begin
        _zz__zz_regVec_0 = regVec_511;
      end
      12'b001000000000 : begin
        _zz__zz_regVec_0 = regVec_512;
      end
      12'b001000000001 : begin
        _zz__zz_regVec_0 = regVec_513;
      end
      12'b001000000010 : begin
        _zz__zz_regVec_0 = regVec_514;
      end
      12'b001000000011 : begin
        _zz__zz_regVec_0 = regVec_515;
      end
      12'b001000000100 : begin
        _zz__zz_regVec_0 = regVec_516;
      end
      12'b001000000101 : begin
        _zz__zz_regVec_0 = regVec_517;
      end
      12'b001000000110 : begin
        _zz__zz_regVec_0 = regVec_518;
      end
      12'b001000000111 : begin
        _zz__zz_regVec_0 = regVec_519;
      end
      12'b001000001000 : begin
        _zz__zz_regVec_0 = regVec_520;
      end
      12'b001000001001 : begin
        _zz__zz_regVec_0 = regVec_521;
      end
      12'b001000001010 : begin
        _zz__zz_regVec_0 = regVec_522;
      end
      12'b001000001011 : begin
        _zz__zz_regVec_0 = regVec_523;
      end
      12'b001000001100 : begin
        _zz__zz_regVec_0 = regVec_524;
      end
      12'b001000001101 : begin
        _zz__zz_regVec_0 = regVec_525;
      end
      12'b001000001110 : begin
        _zz__zz_regVec_0 = regVec_526;
      end
      12'b001000001111 : begin
        _zz__zz_regVec_0 = regVec_527;
      end
      12'b001000010000 : begin
        _zz__zz_regVec_0 = regVec_528;
      end
      12'b001000010001 : begin
        _zz__zz_regVec_0 = regVec_529;
      end
      12'b001000010010 : begin
        _zz__zz_regVec_0 = regVec_530;
      end
      12'b001000010011 : begin
        _zz__zz_regVec_0 = regVec_531;
      end
      12'b001000010100 : begin
        _zz__zz_regVec_0 = regVec_532;
      end
      12'b001000010101 : begin
        _zz__zz_regVec_0 = regVec_533;
      end
      12'b001000010110 : begin
        _zz__zz_regVec_0 = regVec_534;
      end
      12'b001000010111 : begin
        _zz__zz_regVec_0 = regVec_535;
      end
      12'b001000011000 : begin
        _zz__zz_regVec_0 = regVec_536;
      end
      12'b001000011001 : begin
        _zz__zz_regVec_0 = regVec_537;
      end
      12'b001000011010 : begin
        _zz__zz_regVec_0 = regVec_538;
      end
      12'b001000011011 : begin
        _zz__zz_regVec_0 = regVec_539;
      end
      12'b001000011100 : begin
        _zz__zz_regVec_0 = regVec_540;
      end
      12'b001000011101 : begin
        _zz__zz_regVec_0 = regVec_541;
      end
      12'b001000011110 : begin
        _zz__zz_regVec_0 = regVec_542;
      end
      12'b001000011111 : begin
        _zz__zz_regVec_0 = regVec_543;
      end
      12'b001000100000 : begin
        _zz__zz_regVec_0 = regVec_544;
      end
      12'b001000100001 : begin
        _zz__zz_regVec_0 = regVec_545;
      end
      12'b001000100010 : begin
        _zz__zz_regVec_0 = regVec_546;
      end
      12'b001000100011 : begin
        _zz__zz_regVec_0 = regVec_547;
      end
      12'b001000100100 : begin
        _zz__zz_regVec_0 = regVec_548;
      end
      12'b001000100101 : begin
        _zz__zz_regVec_0 = regVec_549;
      end
      12'b001000100110 : begin
        _zz__zz_regVec_0 = regVec_550;
      end
      12'b001000100111 : begin
        _zz__zz_regVec_0 = regVec_551;
      end
      12'b001000101000 : begin
        _zz__zz_regVec_0 = regVec_552;
      end
      12'b001000101001 : begin
        _zz__zz_regVec_0 = regVec_553;
      end
      12'b001000101010 : begin
        _zz__zz_regVec_0 = regVec_554;
      end
      12'b001000101011 : begin
        _zz__zz_regVec_0 = regVec_555;
      end
      12'b001000101100 : begin
        _zz__zz_regVec_0 = regVec_556;
      end
      12'b001000101101 : begin
        _zz__zz_regVec_0 = regVec_557;
      end
      12'b001000101110 : begin
        _zz__zz_regVec_0 = regVec_558;
      end
      12'b001000101111 : begin
        _zz__zz_regVec_0 = regVec_559;
      end
      12'b001000110000 : begin
        _zz__zz_regVec_0 = regVec_560;
      end
      12'b001000110001 : begin
        _zz__zz_regVec_0 = regVec_561;
      end
      12'b001000110010 : begin
        _zz__zz_regVec_0 = regVec_562;
      end
      12'b001000110011 : begin
        _zz__zz_regVec_0 = regVec_563;
      end
      12'b001000110100 : begin
        _zz__zz_regVec_0 = regVec_564;
      end
      12'b001000110101 : begin
        _zz__zz_regVec_0 = regVec_565;
      end
      12'b001000110110 : begin
        _zz__zz_regVec_0 = regVec_566;
      end
      12'b001000110111 : begin
        _zz__zz_regVec_0 = regVec_567;
      end
      12'b001000111000 : begin
        _zz__zz_regVec_0 = regVec_568;
      end
      12'b001000111001 : begin
        _zz__zz_regVec_0 = regVec_569;
      end
      12'b001000111010 : begin
        _zz__zz_regVec_0 = regVec_570;
      end
      12'b001000111011 : begin
        _zz__zz_regVec_0 = regVec_571;
      end
      12'b001000111100 : begin
        _zz__zz_regVec_0 = regVec_572;
      end
      12'b001000111101 : begin
        _zz__zz_regVec_0 = regVec_573;
      end
      12'b001000111110 : begin
        _zz__zz_regVec_0 = regVec_574;
      end
      12'b001000111111 : begin
        _zz__zz_regVec_0 = regVec_575;
      end
      12'b001001000000 : begin
        _zz__zz_regVec_0 = regVec_576;
      end
      12'b001001000001 : begin
        _zz__zz_regVec_0 = regVec_577;
      end
      12'b001001000010 : begin
        _zz__zz_regVec_0 = regVec_578;
      end
      12'b001001000011 : begin
        _zz__zz_regVec_0 = regVec_579;
      end
      12'b001001000100 : begin
        _zz__zz_regVec_0 = regVec_580;
      end
      12'b001001000101 : begin
        _zz__zz_regVec_0 = regVec_581;
      end
      12'b001001000110 : begin
        _zz__zz_regVec_0 = regVec_582;
      end
      12'b001001000111 : begin
        _zz__zz_regVec_0 = regVec_583;
      end
      12'b001001001000 : begin
        _zz__zz_regVec_0 = regVec_584;
      end
      12'b001001001001 : begin
        _zz__zz_regVec_0 = regVec_585;
      end
      12'b001001001010 : begin
        _zz__zz_regVec_0 = regVec_586;
      end
      12'b001001001011 : begin
        _zz__zz_regVec_0 = regVec_587;
      end
      12'b001001001100 : begin
        _zz__zz_regVec_0 = regVec_588;
      end
      12'b001001001101 : begin
        _zz__zz_regVec_0 = regVec_589;
      end
      12'b001001001110 : begin
        _zz__zz_regVec_0 = regVec_590;
      end
      12'b001001001111 : begin
        _zz__zz_regVec_0 = regVec_591;
      end
      12'b001001010000 : begin
        _zz__zz_regVec_0 = regVec_592;
      end
      12'b001001010001 : begin
        _zz__zz_regVec_0 = regVec_593;
      end
      12'b001001010010 : begin
        _zz__zz_regVec_0 = regVec_594;
      end
      12'b001001010011 : begin
        _zz__zz_regVec_0 = regVec_595;
      end
      12'b001001010100 : begin
        _zz__zz_regVec_0 = regVec_596;
      end
      12'b001001010101 : begin
        _zz__zz_regVec_0 = regVec_597;
      end
      12'b001001010110 : begin
        _zz__zz_regVec_0 = regVec_598;
      end
      12'b001001010111 : begin
        _zz__zz_regVec_0 = regVec_599;
      end
      12'b001001011000 : begin
        _zz__zz_regVec_0 = regVec_600;
      end
      12'b001001011001 : begin
        _zz__zz_regVec_0 = regVec_601;
      end
      12'b001001011010 : begin
        _zz__zz_regVec_0 = regVec_602;
      end
      12'b001001011011 : begin
        _zz__zz_regVec_0 = regVec_603;
      end
      12'b001001011100 : begin
        _zz__zz_regVec_0 = regVec_604;
      end
      12'b001001011101 : begin
        _zz__zz_regVec_0 = regVec_605;
      end
      12'b001001011110 : begin
        _zz__zz_regVec_0 = regVec_606;
      end
      12'b001001011111 : begin
        _zz__zz_regVec_0 = regVec_607;
      end
      12'b001001100000 : begin
        _zz__zz_regVec_0 = regVec_608;
      end
      12'b001001100001 : begin
        _zz__zz_regVec_0 = regVec_609;
      end
      12'b001001100010 : begin
        _zz__zz_regVec_0 = regVec_610;
      end
      12'b001001100011 : begin
        _zz__zz_regVec_0 = regVec_611;
      end
      12'b001001100100 : begin
        _zz__zz_regVec_0 = regVec_612;
      end
      12'b001001100101 : begin
        _zz__zz_regVec_0 = regVec_613;
      end
      12'b001001100110 : begin
        _zz__zz_regVec_0 = regVec_614;
      end
      12'b001001100111 : begin
        _zz__zz_regVec_0 = regVec_615;
      end
      12'b001001101000 : begin
        _zz__zz_regVec_0 = regVec_616;
      end
      12'b001001101001 : begin
        _zz__zz_regVec_0 = regVec_617;
      end
      12'b001001101010 : begin
        _zz__zz_regVec_0 = regVec_618;
      end
      12'b001001101011 : begin
        _zz__zz_regVec_0 = regVec_619;
      end
      12'b001001101100 : begin
        _zz__zz_regVec_0 = regVec_620;
      end
      12'b001001101101 : begin
        _zz__zz_regVec_0 = regVec_621;
      end
      12'b001001101110 : begin
        _zz__zz_regVec_0 = regVec_622;
      end
      12'b001001101111 : begin
        _zz__zz_regVec_0 = regVec_623;
      end
      12'b001001110000 : begin
        _zz__zz_regVec_0 = regVec_624;
      end
      12'b001001110001 : begin
        _zz__zz_regVec_0 = regVec_625;
      end
      12'b001001110010 : begin
        _zz__zz_regVec_0 = regVec_626;
      end
      12'b001001110011 : begin
        _zz__zz_regVec_0 = regVec_627;
      end
      12'b001001110100 : begin
        _zz__zz_regVec_0 = regVec_628;
      end
      12'b001001110101 : begin
        _zz__zz_regVec_0 = regVec_629;
      end
      12'b001001110110 : begin
        _zz__zz_regVec_0 = regVec_630;
      end
      12'b001001110111 : begin
        _zz__zz_regVec_0 = regVec_631;
      end
      12'b001001111000 : begin
        _zz__zz_regVec_0 = regVec_632;
      end
      12'b001001111001 : begin
        _zz__zz_regVec_0 = regVec_633;
      end
      12'b001001111010 : begin
        _zz__zz_regVec_0 = regVec_634;
      end
      12'b001001111011 : begin
        _zz__zz_regVec_0 = regVec_635;
      end
      12'b001001111100 : begin
        _zz__zz_regVec_0 = regVec_636;
      end
      12'b001001111101 : begin
        _zz__zz_regVec_0 = regVec_637;
      end
      12'b001001111110 : begin
        _zz__zz_regVec_0 = regVec_638;
      end
      12'b001001111111 : begin
        _zz__zz_regVec_0 = regVec_639;
      end
      12'b001010000000 : begin
        _zz__zz_regVec_0 = regVec_640;
      end
      12'b001010000001 : begin
        _zz__zz_regVec_0 = regVec_641;
      end
      12'b001010000010 : begin
        _zz__zz_regVec_0 = regVec_642;
      end
      12'b001010000011 : begin
        _zz__zz_regVec_0 = regVec_643;
      end
      12'b001010000100 : begin
        _zz__zz_regVec_0 = regVec_644;
      end
      12'b001010000101 : begin
        _zz__zz_regVec_0 = regVec_645;
      end
      12'b001010000110 : begin
        _zz__zz_regVec_0 = regVec_646;
      end
      12'b001010000111 : begin
        _zz__zz_regVec_0 = regVec_647;
      end
      12'b001010001000 : begin
        _zz__zz_regVec_0 = regVec_648;
      end
      12'b001010001001 : begin
        _zz__zz_regVec_0 = regVec_649;
      end
      12'b001010001010 : begin
        _zz__zz_regVec_0 = regVec_650;
      end
      12'b001010001011 : begin
        _zz__zz_regVec_0 = regVec_651;
      end
      12'b001010001100 : begin
        _zz__zz_regVec_0 = regVec_652;
      end
      12'b001010001101 : begin
        _zz__zz_regVec_0 = regVec_653;
      end
      12'b001010001110 : begin
        _zz__zz_regVec_0 = regVec_654;
      end
      12'b001010001111 : begin
        _zz__zz_regVec_0 = regVec_655;
      end
      12'b001010010000 : begin
        _zz__zz_regVec_0 = regVec_656;
      end
      12'b001010010001 : begin
        _zz__zz_regVec_0 = regVec_657;
      end
      12'b001010010010 : begin
        _zz__zz_regVec_0 = regVec_658;
      end
      12'b001010010011 : begin
        _zz__zz_regVec_0 = regVec_659;
      end
      12'b001010010100 : begin
        _zz__zz_regVec_0 = regVec_660;
      end
      12'b001010010101 : begin
        _zz__zz_regVec_0 = regVec_661;
      end
      12'b001010010110 : begin
        _zz__zz_regVec_0 = regVec_662;
      end
      12'b001010010111 : begin
        _zz__zz_regVec_0 = regVec_663;
      end
      12'b001010011000 : begin
        _zz__zz_regVec_0 = regVec_664;
      end
      12'b001010011001 : begin
        _zz__zz_regVec_0 = regVec_665;
      end
      12'b001010011010 : begin
        _zz__zz_regVec_0 = regVec_666;
      end
      12'b001010011011 : begin
        _zz__zz_regVec_0 = regVec_667;
      end
      12'b001010011100 : begin
        _zz__zz_regVec_0 = regVec_668;
      end
      12'b001010011101 : begin
        _zz__zz_regVec_0 = regVec_669;
      end
      12'b001010011110 : begin
        _zz__zz_regVec_0 = regVec_670;
      end
      12'b001010011111 : begin
        _zz__zz_regVec_0 = regVec_671;
      end
      12'b001010100000 : begin
        _zz__zz_regVec_0 = regVec_672;
      end
      12'b001010100001 : begin
        _zz__zz_regVec_0 = regVec_673;
      end
      12'b001010100010 : begin
        _zz__zz_regVec_0 = regVec_674;
      end
      12'b001010100011 : begin
        _zz__zz_regVec_0 = regVec_675;
      end
      12'b001010100100 : begin
        _zz__zz_regVec_0 = regVec_676;
      end
      12'b001010100101 : begin
        _zz__zz_regVec_0 = regVec_677;
      end
      12'b001010100110 : begin
        _zz__zz_regVec_0 = regVec_678;
      end
      12'b001010100111 : begin
        _zz__zz_regVec_0 = regVec_679;
      end
      12'b001010101000 : begin
        _zz__zz_regVec_0 = regVec_680;
      end
      12'b001010101001 : begin
        _zz__zz_regVec_0 = regVec_681;
      end
      12'b001010101010 : begin
        _zz__zz_regVec_0 = regVec_682;
      end
      12'b001010101011 : begin
        _zz__zz_regVec_0 = regVec_683;
      end
      12'b001010101100 : begin
        _zz__zz_regVec_0 = regVec_684;
      end
      12'b001010101101 : begin
        _zz__zz_regVec_0 = regVec_685;
      end
      12'b001010101110 : begin
        _zz__zz_regVec_0 = regVec_686;
      end
      12'b001010101111 : begin
        _zz__zz_regVec_0 = regVec_687;
      end
      12'b001010110000 : begin
        _zz__zz_regVec_0 = regVec_688;
      end
      12'b001010110001 : begin
        _zz__zz_regVec_0 = regVec_689;
      end
      12'b001010110010 : begin
        _zz__zz_regVec_0 = regVec_690;
      end
      12'b001010110011 : begin
        _zz__zz_regVec_0 = regVec_691;
      end
      12'b001010110100 : begin
        _zz__zz_regVec_0 = regVec_692;
      end
      12'b001010110101 : begin
        _zz__zz_regVec_0 = regVec_693;
      end
      12'b001010110110 : begin
        _zz__zz_regVec_0 = regVec_694;
      end
      12'b001010110111 : begin
        _zz__zz_regVec_0 = regVec_695;
      end
      12'b001010111000 : begin
        _zz__zz_regVec_0 = regVec_696;
      end
      12'b001010111001 : begin
        _zz__zz_regVec_0 = regVec_697;
      end
      12'b001010111010 : begin
        _zz__zz_regVec_0 = regVec_698;
      end
      12'b001010111011 : begin
        _zz__zz_regVec_0 = regVec_699;
      end
      12'b001010111100 : begin
        _zz__zz_regVec_0 = regVec_700;
      end
      12'b001010111101 : begin
        _zz__zz_regVec_0 = regVec_701;
      end
      12'b001010111110 : begin
        _zz__zz_regVec_0 = regVec_702;
      end
      12'b001010111111 : begin
        _zz__zz_regVec_0 = regVec_703;
      end
      12'b001011000000 : begin
        _zz__zz_regVec_0 = regVec_704;
      end
      12'b001011000001 : begin
        _zz__zz_regVec_0 = regVec_705;
      end
      12'b001011000010 : begin
        _zz__zz_regVec_0 = regVec_706;
      end
      12'b001011000011 : begin
        _zz__zz_regVec_0 = regVec_707;
      end
      12'b001011000100 : begin
        _zz__zz_regVec_0 = regVec_708;
      end
      12'b001011000101 : begin
        _zz__zz_regVec_0 = regVec_709;
      end
      12'b001011000110 : begin
        _zz__zz_regVec_0 = regVec_710;
      end
      12'b001011000111 : begin
        _zz__zz_regVec_0 = regVec_711;
      end
      12'b001011001000 : begin
        _zz__zz_regVec_0 = regVec_712;
      end
      12'b001011001001 : begin
        _zz__zz_regVec_0 = regVec_713;
      end
      12'b001011001010 : begin
        _zz__zz_regVec_0 = regVec_714;
      end
      12'b001011001011 : begin
        _zz__zz_regVec_0 = regVec_715;
      end
      12'b001011001100 : begin
        _zz__zz_regVec_0 = regVec_716;
      end
      12'b001011001101 : begin
        _zz__zz_regVec_0 = regVec_717;
      end
      12'b001011001110 : begin
        _zz__zz_regVec_0 = regVec_718;
      end
      12'b001011001111 : begin
        _zz__zz_regVec_0 = regVec_719;
      end
      12'b001011010000 : begin
        _zz__zz_regVec_0 = regVec_720;
      end
      12'b001011010001 : begin
        _zz__zz_regVec_0 = regVec_721;
      end
      12'b001011010010 : begin
        _zz__zz_regVec_0 = regVec_722;
      end
      12'b001011010011 : begin
        _zz__zz_regVec_0 = regVec_723;
      end
      12'b001011010100 : begin
        _zz__zz_regVec_0 = regVec_724;
      end
      12'b001011010101 : begin
        _zz__zz_regVec_0 = regVec_725;
      end
      12'b001011010110 : begin
        _zz__zz_regVec_0 = regVec_726;
      end
      12'b001011010111 : begin
        _zz__zz_regVec_0 = regVec_727;
      end
      12'b001011011000 : begin
        _zz__zz_regVec_0 = regVec_728;
      end
      12'b001011011001 : begin
        _zz__zz_regVec_0 = regVec_729;
      end
      12'b001011011010 : begin
        _zz__zz_regVec_0 = regVec_730;
      end
      12'b001011011011 : begin
        _zz__zz_regVec_0 = regVec_731;
      end
      12'b001011011100 : begin
        _zz__zz_regVec_0 = regVec_732;
      end
      12'b001011011101 : begin
        _zz__zz_regVec_0 = regVec_733;
      end
      12'b001011011110 : begin
        _zz__zz_regVec_0 = regVec_734;
      end
      12'b001011011111 : begin
        _zz__zz_regVec_0 = regVec_735;
      end
      12'b001011100000 : begin
        _zz__zz_regVec_0 = regVec_736;
      end
      12'b001011100001 : begin
        _zz__zz_regVec_0 = regVec_737;
      end
      12'b001011100010 : begin
        _zz__zz_regVec_0 = regVec_738;
      end
      12'b001011100011 : begin
        _zz__zz_regVec_0 = regVec_739;
      end
      12'b001011100100 : begin
        _zz__zz_regVec_0 = regVec_740;
      end
      12'b001011100101 : begin
        _zz__zz_regVec_0 = regVec_741;
      end
      12'b001011100110 : begin
        _zz__zz_regVec_0 = regVec_742;
      end
      12'b001011100111 : begin
        _zz__zz_regVec_0 = regVec_743;
      end
      12'b001011101000 : begin
        _zz__zz_regVec_0 = regVec_744;
      end
      12'b001011101001 : begin
        _zz__zz_regVec_0 = regVec_745;
      end
      12'b001011101010 : begin
        _zz__zz_regVec_0 = regVec_746;
      end
      12'b001011101011 : begin
        _zz__zz_regVec_0 = regVec_747;
      end
      12'b001011101100 : begin
        _zz__zz_regVec_0 = regVec_748;
      end
      12'b001011101101 : begin
        _zz__zz_regVec_0 = regVec_749;
      end
      12'b001011101110 : begin
        _zz__zz_regVec_0 = regVec_750;
      end
      12'b001011101111 : begin
        _zz__zz_regVec_0 = regVec_751;
      end
      12'b001011110000 : begin
        _zz__zz_regVec_0 = regVec_752;
      end
      12'b001011110001 : begin
        _zz__zz_regVec_0 = regVec_753;
      end
      12'b001011110010 : begin
        _zz__zz_regVec_0 = regVec_754;
      end
      12'b001011110011 : begin
        _zz__zz_regVec_0 = regVec_755;
      end
      12'b001011110100 : begin
        _zz__zz_regVec_0 = regVec_756;
      end
      12'b001011110101 : begin
        _zz__zz_regVec_0 = regVec_757;
      end
      12'b001011110110 : begin
        _zz__zz_regVec_0 = regVec_758;
      end
      12'b001011110111 : begin
        _zz__zz_regVec_0 = regVec_759;
      end
      12'b001011111000 : begin
        _zz__zz_regVec_0 = regVec_760;
      end
      12'b001011111001 : begin
        _zz__zz_regVec_0 = regVec_761;
      end
      12'b001011111010 : begin
        _zz__zz_regVec_0 = regVec_762;
      end
      12'b001011111011 : begin
        _zz__zz_regVec_0 = regVec_763;
      end
      12'b001011111100 : begin
        _zz__zz_regVec_0 = regVec_764;
      end
      12'b001011111101 : begin
        _zz__zz_regVec_0 = regVec_765;
      end
      12'b001011111110 : begin
        _zz__zz_regVec_0 = regVec_766;
      end
      12'b001011111111 : begin
        _zz__zz_regVec_0 = regVec_767;
      end
      12'b001100000000 : begin
        _zz__zz_regVec_0 = regVec_768;
      end
      12'b001100000001 : begin
        _zz__zz_regVec_0 = regVec_769;
      end
      12'b001100000010 : begin
        _zz__zz_regVec_0 = regVec_770;
      end
      12'b001100000011 : begin
        _zz__zz_regVec_0 = regVec_771;
      end
      12'b001100000100 : begin
        _zz__zz_regVec_0 = regVec_772;
      end
      12'b001100000101 : begin
        _zz__zz_regVec_0 = regVec_773;
      end
      12'b001100000110 : begin
        _zz__zz_regVec_0 = regVec_774;
      end
      12'b001100000111 : begin
        _zz__zz_regVec_0 = regVec_775;
      end
      12'b001100001000 : begin
        _zz__zz_regVec_0 = regVec_776;
      end
      12'b001100001001 : begin
        _zz__zz_regVec_0 = regVec_777;
      end
      12'b001100001010 : begin
        _zz__zz_regVec_0 = regVec_778;
      end
      12'b001100001011 : begin
        _zz__zz_regVec_0 = regVec_779;
      end
      12'b001100001100 : begin
        _zz__zz_regVec_0 = regVec_780;
      end
      12'b001100001101 : begin
        _zz__zz_regVec_0 = regVec_781;
      end
      12'b001100001110 : begin
        _zz__zz_regVec_0 = regVec_782;
      end
      12'b001100001111 : begin
        _zz__zz_regVec_0 = regVec_783;
      end
      12'b001100010000 : begin
        _zz__zz_regVec_0 = regVec_784;
      end
      12'b001100010001 : begin
        _zz__zz_regVec_0 = regVec_785;
      end
      12'b001100010010 : begin
        _zz__zz_regVec_0 = regVec_786;
      end
      12'b001100010011 : begin
        _zz__zz_regVec_0 = regVec_787;
      end
      12'b001100010100 : begin
        _zz__zz_regVec_0 = regVec_788;
      end
      12'b001100010101 : begin
        _zz__zz_regVec_0 = regVec_789;
      end
      12'b001100010110 : begin
        _zz__zz_regVec_0 = regVec_790;
      end
      12'b001100010111 : begin
        _zz__zz_regVec_0 = regVec_791;
      end
      12'b001100011000 : begin
        _zz__zz_regVec_0 = regVec_792;
      end
      12'b001100011001 : begin
        _zz__zz_regVec_0 = regVec_793;
      end
      12'b001100011010 : begin
        _zz__zz_regVec_0 = regVec_794;
      end
      12'b001100011011 : begin
        _zz__zz_regVec_0 = regVec_795;
      end
      12'b001100011100 : begin
        _zz__zz_regVec_0 = regVec_796;
      end
      12'b001100011101 : begin
        _zz__zz_regVec_0 = regVec_797;
      end
      12'b001100011110 : begin
        _zz__zz_regVec_0 = regVec_798;
      end
      12'b001100011111 : begin
        _zz__zz_regVec_0 = regVec_799;
      end
      12'b001100100000 : begin
        _zz__zz_regVec_0 = regVec_800;
      end
      12'b001100100001 : begin
        _zz__zz_regVec_0 = regVec_801;
      end
      12'b001100100010 : begin
        _zz__zz_regVec_0 = regVec_802;
      end
      12'b001100100011 : begin
        _zz__zz_regVec_0 = regVec_803;
      end
      12'b001100100100 : begin
        _zz__zz_regVec_0 = regVec_804;
      end
      12'b001100100101 : begin
        _zz__zz_regVec_0 = regVec_805;
      end
      12'b001100100110 : begin
        _zz__zz_regVec_0 = regVec_806;
      end
      12'b001100100111 : begin
        _zz__zz_regVec_0 = regVec_807;
      end
      12'b001100101000 : begin
        _zz__zz_regVec_0 = regVec_808;
      end
      12'b001100101001 : begin
        _zz__zz_regVec_0 = regVec_809;
      end
      12'b001100101010 : begin
        _zz__zz_regVec_0 = regVec_810;
      end
      12'b001100101011 : begin
        _zz__zz_regVec_0 = regVec_811;
      end
      12'b001100101100 : begin
        _zz__zz_regVec_0 = regVec_812;
      end
      12'b001100101101 : begin
        _zz__zz_regVec_0 = regVec_813;
      end
      12'b001100101110 : begin
        _zz__zz_regVec_0 = regVec_814;
      end
      12'b001100101111 : begin
        _zz__zz_regVec_0 = regVec_815;
      end
      12'b001100110000 : begin
        _zz__zz_regVec_0 = regVec_816;
      end
      12'b001100110001 : begin
        _zz__zz_regVec_0 = regVec_817;
      end
      12'b001100110010 : begin
        _zz__zz_regVec_0 = regVec_818;
      end
      12'b001100110011 : begin
        _zz__zz_regVec_0 = regVec_819;
      end
      12'b001100110100 : begin
        _zz__zz_regVec_0 = regVec_820;
      end
      12'b001100110101 : begin
        _zz__zz_regVec_0 = regVec_821;
      end
      12'b001100110110 : begin
        _zz__zz_regVec_0 = regVec_822;
      end
      12'b001100110111 : begin
        _zz__zz_regVec_0 = regVec_823;
      end
      12'b001100111000 : begin
        _zz__zz_regVec_0 = regVec_824;
      end
      12'b001100111001 : begin
        _zz__zz_regVec_0 = regVec_825;
      end
      12'b001100111010 : begin
        _zz__zz_regVec_0 = regVec_826;
      end
      12'b001100111011 : begin
        _zz__zz_regVec_0 = regVec_827;
      end
      12'b001100111100 : begin
        _zz__zz_regVec_0 = regVec_828;
      end
      12'b001100111101 : begin
        _zz__zz_regVec_0 = regVec_829;
      end
      12'b001100111110 : begin
        _zz__zz_regVec_0 = regVec_830;
      end
      12'b001100111111 : begin
        _zz__zz_regVec_0 = regVec_831;
      end
      12'b001101000000 : begin
        _zz__zz_regVec_0 = regVec_832;
      end
      12'b001101000001 : begin
        _zz__zz_regVec_0 = regVec_833;
      end
      12'b001101000010 : begin
        _zz__zz_regVec_0 = regVec_834;
      end
      12'b001101000011 : begin
        _zz__zz_regVec_0 = regVec_835;
      end
      12'b001101000100 : begin
        _zz__zz_regVec_0 = regVec_836;
      end
      12'b001101000101 : begin
        _zz__zz_regVec_0 = regVec_837;
      end
      12'b001101000110 : begin
        _zz__zz_regVec_0 = regVec_838;
      end
      12'b001101000111 : begin
        _zz__zz_regVec_0 = regVec_839;
      end
      12'b001101001000 : begin
        _zz__zz_regVec_0 = regVec_840;
      end
      12'b001101001001 : begin
        _zz__zz_regVec_0 = regVec_841;
      end
      12'b001101001010 : begin
        _zz__zz_regVec_0 = regVec_842;
      end
      12'b001101001011 : begin
        _zz__zz_regVec_0 = regVec_843;
      end
      12'b001101001100 : begin
        _zz__zz_regVec_0 = regVec_844;
      end
      12'b001101001101 : begin
        _zz__zz_regVec_0 = regVec_845;
      end
      12'b001101001110 : begin
        _zz__zz_regVec_0 = regVec_846;
      end
      12'b001101001111 : begin
        _zz__zz_regVec_0 = regVec_847;
      end
      12'b001101010000 : begin
        _zz__zz_regVec_0 = regVec_848;
      end
      12'b001101010001 : begin
        _zz__zz_regVec_0 = regVec_849;
      end
      12'b001101010010 : begin
        _zz__zz_regVec_0 = regVec_850;
      end
      12'b001101010011 : begin
        _zz__zz_regVec_0 = regVec_851;
      end
      12'b001101010100 : begin
        _zz__zz_regVec_0 = regVec_852;
      end
      12'b001101010101 : begin
        _zz__zz_regVec_0 = regVec_853;
      end
      12'b001101010110 : begin
        _zz__zz_regVec_0 = regVec_854;
      end
      12'b001101010111 : begin
        _zz__zz_regVec_0 = regVec_855;
      end
      12'b001101011000 : begin
        _zz__zz_regVec_0 = regVec_856;
      end
      12'b001101011001 : begin
        _zz__zz_regVec_0 = regVec_857;
      end
      12'b001101011010 : begin
        _zz__zz_regVec_0 = regVec_858;
      end
      12'b001101011011 : begin
        _zz__zz_regVec_0 = regVec_859;
      end
      12'b001101011100 : begin
        _zz__zz_regVec_0 = regVec_860;
      end
      12'b001101011101 : begin
        _zz__zz_regVec_0 = regVec_861;
      end
      12'b001101011110 : begin
        _zz__zz_regVec_0 = regVec_862;
      end
      12'b001101011111 : begin
        _zz__zz_regVec_0 = regVec_863;
      end
      12'b001101100000 : begin
        _zz__zz_regVec_0 = regVec_864;
      end
      12'b001101100001 : begin
        _zz__zz_regVec_0 = regVec_865;
      end
      12'b001101100010 : begin
        _zz__zz_regVec_0 = regVec_866;
      end
      12'b001101100011 : begin
        _zz__zz_regVec_0 = regVec_867;
      end
      12'b001101100100 : begin
        _zz__zz_regVec_0 = regVec_868;
      end
      12'b001101100101 : begin
        _zz__zz_regVec_0 = regVec_869;
      end
      12'b001101100110 : begin
        _zz__zz_regVec_0 = regVec_870;
      end
      12'b001101100111 : begin
        _zz__zz_regVec_0 = regVec_871;
      end
      12'b001101101000 : begin
        _zz__zz_regVec_0 = regVec_872;
      end
      12'b001101101001 : begin
        _zz__zz_regVec_0 = regVec_873;
      end
      12'b001101101010 : begin
        _zz__zz_regVec_0 = regVec_874;
      end
      12'b001101101011 : begin
        _zz__zz_regVec_0 = regVec_875;
      end
      12'b001101101100 : begin
        _zz__zz_regVec_0 = regVec_876;
      end
      12'b001101101101 : begin
        _zz__zz_regVec_0 = regVec_877;
      end
      12'b001101101110 : begin
        _zz__zz_regVec_0 = regVec_878;
      end
      12'b001101101111 : begin
        _zz__zz_regVec_0 = regVec_879;
      end
      12'b001101110000 : begin
        _zz__zz_regVec_0 = regVec_880;
      end
      12'b001101110001 : begin
        _zz__zz_regVec_0 = regVec_881;
      end
      12'b001101110010 : begin
        _zz__zz_regVec_0 = regVec_882;
      end
      12'b001101110011 : begin
        _zz__zz_regVec_0 = regVec_883;
      end
      12'b001101110100 : begin
        _zz__zz_regVec_0 = regVec_884;
      end
      12'b001101110101 : begin
        _zz__zz_regVec_0 = regVec_885;
      end
      12'b001101110110 : begin
        _zz__zz_regVec_0 = regVec_886;
      end
      12'b001101110111 : begin
        _zz__zz_regVec_0 = regVec_887;
      end
      12'b001101111000 : begin
        _zz__zz_regVec_0 = regVec_888;
      end
      12'b001101111001 : begin
        _zz__zz_regVec_0 = regVec_889;
      end
      12'b001101111010 : begin
        _zz__zz_regVec_0 = regVec_890;
      end
      12'b001101111011 : begin
        _zz__zz_regVec_0 = regVec_891;
      end
      12'b001101111100 : begin
        _zz__zz_regVec_0 = regVec_892;
      end
      12'b001101111101 : begin
        _zz__zz_regVec_0 = regVec_893;
      end
      12'b001101111110 : begin
        _zz__zz_regVec_0 = regVec_894;
      end
      12'b001101111111 : begin
        _zz__zz_regVec_0 = regVec_895;
      end
      12'b001110000000 : begin
        _zz__zz_regVec_0 = regVec_896;
      end
      12'b001110000001 : begin
        _zz__zz_regVec_0 = regVec_897;
      end
      12'b001110000010 : begin
        _zz__zz_regVec_0 = regVec_898;
      end
      12'b001110000011 : begin
        _zz__zz_regVec_0 = regVec_899;
      end
      12'b001110000100 : begin
        _zz__zz_regVec_0 = regVec_900;
      end
      12'b001110000101 : begin
        _zz__zz_regVec_0 = regVec_901;
      end
      12'b001110000110 : begin
        _zz__zz_regVec_0 = regVec_902;
      end
      12'b001110000111 : begin
        _zz__zz_regVec_0 = regVec_903;
      end
      12'b001110001000 : begin
        _zz__zz_regVec_0 = regVec_904;
      end
      12'b001110001001 : begin
        _zz__zz_regVec_0 = regVec_905;
      end
      12'b001110001010 : begin
        _zz__zz_regVec_0 = regVec_906;
      end
      12'b001110001011 : begin
        _zz__zz_regVec_0 = regVec_907;
      end
      12'b001110001100 : begin
        _zz__zz_regVec_0 = regVec_908;
      end
      12'b001110001101 : begin
        _zz__zz_regVec_0 = regVec_909;
      end
      12'b001110001110 : begin
        _zz__zz_regVec_0 = regVec_910;
      end
      12'b001110001111 : begin
        _zz__zz_regVec_0 = regVec_911;
      end
      12'b001110010000 : begin
        _zz__zz_regVec_0 = regVec_912;
      end
      12'b001110010001 : begin
        _zz__zz_regVec_0 = regVec_913;
      end
      12'b001110010010 : begin
        _zz__zz_regVec_0 = regVec_914;
      end
      12'b001110010011 : begin
        _zz__zz_regVec_0 = regVec_915;
      end
      12'b001110010100 : begin
        _zz__zz_regVec_0 = regVec_916;
      end
      12'b001110010101 : begin
        _zz__zz_regVec_0 = regVec_917;
      end
      12'b001110010110 : begin
        _zz__zz_regVec_0 = regVec_918;
      end
      12'b001110010111 : begin
        _zz__zz_regVec_0 = regVec_919;
      end
      12'b001110011000 : begin
        _zz__zz_regVec_0 = regVec_920;
      end
      12'b001110011001 : begin
        _zz__zz_regVec_0 = regVec_921;
      end
      12'b001110011010 : begin
        _zz__zz_regVec_0 = regVec_922;
      end
      12'b001110011011 : begin
        _zz__zz_regVec_0 = regVec_923;
      end
      12'b001110011100 : begin
        _zz__zz_regVec_0 = regVec_924;
      end
      12'b001110011101 : begin
        _zz__zz_regVec_0 = regVec_925;
      end
      12'b001110011110 : begin
        _zz__zz_regVec_0 = regVec_926;
      end
      12'b001110011111 : begin
        _zz__zz_regVec_0 = regVec_927;
      end
      12'b001110100000 : begin
        _zz__zz_regVec_0 = regVec_928;
      end
      12'b001110100001 : begin
        _zz__zz_regVec_0 = regVec_929;
      end
      12'b001110100010 : begin
        _zz__zz_regVec_0 = regVec_930;
      end
      12'b001110100011 : begin
        _zz__zz_regVec_0 = regVec_931;
      end
      12'b001110100100 : begin
        _zz__zz_regVec_0 = regVec_932;
      end
      12'b001110100101 : begin
        _zz__zz_regVec_0 = regVec_933;
      end
      12'b001110100110 : begin
        _zz__zz_regVec_0 = regVec_934;
      end
      12'b001110100111 : begin
        _zz__zz_regVec_0 = regVec_935;
      end
      12'b001110101000 : begin
        _zz__zz_regVec_0 = regVec_936;
      end
      12'b001110101001 : begin
        _zz__zz_regVec_0 = regVec_937;
      end
      12'b001110101010 : begin
        _zz__zz_regVec_0 = regVec_938;
      end
      12'b001110101011 : begin
        _zz__zz_regVec_0 = regVec_939;
      end
      12'b001110101100 : begin
        _zz__zz_regVec_0 = regVec_940;
      end
      12'b001110101101 : begin
        _zz__zz_regVec_0 = regVec_941;
      end
      12'b001110101110 : begin
        _zz__zz_regVec_0 = regVec_942;
      end
      12'b001110101111 : begin
        _zz__zz_regVec_0 = regVec_943;
      end
      12'b001110110000 : begin
        _zz__zz_regVec_0 = regVec_944;
      end
      12'b001110110001 : begin
        _zz__zz_regVec_0 = regVec_945;
      end
      12'b001110110010 : begin
        _zz__zz_regVec_0 = regVec_946;
      end
      12'b001110110011 : begin
        _zz__zz_regVec_0 = regVec_947;
      end
      12'b001110110100 : begin
        _zz__zz_regVec_0 = regVec_948;
      end
      12'b001110110101 : begin
        _zz__zz_regVec_0 = regVec_949;
      end
      12'b001110110110 : begin
        _zz__zz_regVec_0 = regVec_950;
      end
      12'b001110110111 : begin
        _zz__zz_regVec_0 = regVec_951;
      end
      12'b001110111000 : begin
        _zz__zz_regVec_0 = regVec_952;
      end
      12'b001110111001 : begin
        _zz__zz_regVec_0 = regVec_953;
      end
      12'b001110111010 : begin
        _zz__zz_regVec_0 = regVec_954;
      end
      12'b001110111011 : begin
        _zz__zz_regVec_0 = regVec_955;
      end
      12'b001110111100 : begin
        _zz__zz_regVec_0 = regVec_956;
      end
      12'b001110111101 : begin
        _zz__zz_regVec_0 = regVec_957;
      end
      12'b001110111110 : begin
        _zz__zz_regVec_0 = regVec_958;
      end
      12'b001110111111 : begin
        _zz__zz_regVec_0 = regVec_959;
      end
      12'b001111000000 : begin
        _zz__zz_regVec_0 = regVec_960;
      end
      12'b001111000001 : begin
        _zz__zz_regVec_0 = regVec_961;
      end
      12'b001111000010 : begin
        _zz__zz_regVec_0 = regVec_962;
      end
      12'b001111000011 : begin
        _zz__zz_regVec_0 = regVec_963;
      end
      12'b001111000100 : begin
        _zz__zz_regVec_0 = regVec_964;
      end
      12'b001111000101 : begin
        _zz__zz_regVec_0 = regVec_965;
      end
      12'b001111000110 : begin
        _zz__zz_regVec_0 = regVec_966;
      end
      12'b001111000111 : begin
        _zz__zz_regVec_0 = regVec_967;
      end
      12'b001111001000 : begin
        _zz__zz_regVec_0 = regVec_968;
      end
      12'b001111001001 : begin
        _zz__zz_regVec_0 = regVec_969;
      end
      12'b001111001010 : begin
        _zz__zz_regVec_0 = regVec_970;
      end
      12'b001111001011 : begin
        _zz__zz_regVec_0 = regVec_971;
      end
      12'b001111001100 : begin
        _zz__zz_regVec_0 = regVec_972;
      end
      12'b001111001101 : begin
        _zz__zz_regVec_0 = regVec_973;
      end
      12'b001111001110 : begin
        _zz__zz_regVec_0 = regVec_974;
      end
      12'b001111001111 : begin
        _zz__zz_regVec_0 = regVec_975;
      end
      12'b001111010000 : begin
        _zz__zz_regVec_0 = regVec_976;
      end
      12'b001111010001 : begin
        _zz__zz_regVec_0 = regVec_977;
      end
      12'b001111010010 : begin
        _zz__zz_regVec_0 = regVec_978;
      end
      12'b001111010011 : begin
        _zz__zz_regVec_0 = regVec_979;
      end
      12'b001111010100 : begin
        _zz__zz_regVec_0 = regVec_980;
      end
      12'b001111010101 : begin
        _zz__zz_regVec_0 = regVec_981;
      end
      12'b001111010110 : begin
        _zz__zz_regVec_0 = regVec_982;
      end
      12'b001111010111 : begin
        _zz__zz_regVec_0 = regVec_983;
      end
      12'b001111011000 : begin
        _zz__zz_regVec_0 = regVec_984;
      end
      12'b001111011001 : begin
        _zz__zz_regVec_0 = regVec_985;
      end
      12'b001111011010 : begin
        _zz__zz_regVec_0 = regVec_986;
      end
      12'b001111011011 : begin
        _zz__zz_regVec_0 = regVec_987;
      end
      12'b001111011100 : begin
        _zz__zz_regVec_0 = regVec_988;
      end
      12'b001111011101 : begin
        _zz__zz_regVec_0 = regVec_989;
      end
      12'b001111011110 : begin
        _zz__zz_regVec_0 = regVec_990;
      end
      12'b001111011111 : begin
        _zz__zz_regVec_0 = regVec_991;
      end
      12'b001111100000 : begin
        _zz__zz_regVec_0 = regVec_992;
      end
      12'b001111100001 : begin
        _zz__zz_regVec_0 = regVec_993;
      end
      12'b001111100010 : begin
        _zz__zz_regVec_0 = regVec_994;
      end
      12'b001111100011 : begin
        _zz__zz_regVec_0 = regVec_995;
      end
      12'b001111100100 : begin
        _zz__zz_regVec_0 = regVec_996;
      end
      12'b001111100101 : begin
        _zz__zz_regVec_0 = regVec_997;
      end
      12'b001111100110 : begin
        _zz__zz_regVec_0 = regVec_998;
      end
      12'b001111100111 : begin
        _zz__zz_regVec_0 = regVec_999;
      end
      12'b001111101000 : begin
        _zz__zz_regVec_0 = regVec_1000;
      end
      12'b001111101001 : begin
        _zz__zz_regVec_0 = regVec_1001;
      end
      12'b001111101010 : begin
        _zz__zz_regVec_0 = regVec_1002;
      end
      12'b001111101011 : begin
        _zz__zz_regVec_0 = regVec_1003;
      end
      12'b001111101100 : begin
        _zz__zz_regVec_0 = regVec_1004;
      end
      12'b001111101101 : begin
        _zz__zz_regVec_0 = regVec_1005;
      end
      12'b001111101110 : begin
        _zz__zz_regVec_0 = regVec_1006;
      end
      12'b001111101111 : begin
        _zz__zz_regVec_0 = regVec_1007;
      end
      12'b001111110000 : begin
        _zz__zz_regVec_0 = regVec_1008;
      end
      12'b001111110001 : begin
        _zz__zz_regVec_0 = regVec_1009;
      end
      12'b001111110010 : begin
        _zz__zz_regVec_0 = regVec_1010;
      end
      12'b001111110011 : begin
        _zz__zz_regVec_0 = regVec_1011;
      end
      12'b001111110100 : begin
        _zz__zz_regVec_0 = regVec_1012;
      end
      12'b001111110101 : begin
        _zz__zz_regVec_0 = regVec_1013;
      end
      12'b001111110110 : begin
        _zz__zz_regVec_0 = regVec_1014;
      end
      12'b001111110111 : begin
        _zz__zz_regVec_0 = regVec_1015;
      end
      12'b001111111000 : begin
        _zz__zz_regVec_0 = regVec_1016;
      end
      12'b001111111001 : begin
        _zz__zz_regVec_0 = regVec_1017;
      end
      12'b001111111010 : begin
        _zz__zz_regVec_0 = regVec_1018;
      end
      12'b001111111011 : begin
        _zz__zz_regVec_0 = regVec_1019;
      end
      12'b001111111100 : begin
        _zz__zz_regVec_0 = regVec_1020;
      end
      12'b001111111101 : begin
        _zz__zz_regVec_0 = regVec_1021;
      end
      12'b001111111110 : begin
        _zz__zz_regVec_0 = regVec_1022;
      end
      12'b001111111111 : begin
        _zz__zz_regVec_0 = regVec_1023;
      end
      12'b010000000000 : begin
        _zz__zz_regVec_0 = regVec_1024;
      end
      12'b010000000001 : begin
        _zz__zz_regVec_0 = regVec_1025;
      end
      12'b010000000010 : begin
        _zz__zz_regVec_0 = regVec_1026;
      end
      12'b010000000011 : begin
        _zz__zz_regVec_0 = regVec_1027;
      end
      12'b010000000100 : begin
        _zz__zz_regVec_0 = regVec_1028;
      end
      12'b010000000101 : begin
        _zz__zz_regVec_0 = regVec_1029;
      end
      12'b010000000110 : begin
        _zz__zz_regVec_0 = regVec_1030;
      end
      12'b010000000111 : begin
        _zz__zz_regVec_0 = regVec_1031;
      end
      12'b010000001000 : begin
        _zz__zz_regVec_0 = regVec_1032;
      end
      12'b010000001001 : begin
        _zz__zz_regVec_0 = regVec_1033;
      end
      12'b010000001010 : begin
        _zz__zz_regVec_0 = regVec_1034;
      end
      12'b010000001011 : begin
        _zz__zz_regVec_0 = regVec_1035;
      end
      12'b010000001100 : begin
        _zz__zz_regVec_0 = regVec_1036;
      end
      12'b010000001101 : begin
        _zz__zz_regVec_0 = regVec_1037;
      end
      12'b010000001110 : begin
        _zz__zz_regVec_0 = regVec_1038;
      end
      12'b010000001111 : begin
        _zz__zz_regVec_0 = regVec_1039;
      end
      12'b010000010000 : begin
        _zz__zz_regVec_0 = regVec_1040;
      end
      12'b010000010001 : begin
        _zz__zz_regVec_0 = regVec_1041;
      end
      12'b010000010010 : begin
        _zz__zz_regVec_0 = regVec_1042;
      end
      12'b010000010011 : begin
        _zz__zz_regVec_0 = regVec_1043;
      end
      12'b010000010100 : begin
        _zz__zz_regVec_0 = regVec_1044;
      end
      12'b010000010101 : begin
        _zz__zz_regVec_0 = regVec_1045;
      end
      12'b010000010110 : begin
        _zz__zz_regVec_0 = regVec_1046;
      end
      12'b010000010111 : begin
        _zz__zz_regVec_0 = regVec_1047;
      end
      12'b010000011000 : begin
        _zz__zz_regVec_0 = regVec_1048;
      end
      12'b010000011001 : begin
        _zz__zz_regVec_0 = regVec_1049;
      end
      12'b010000011010 : begin
        _zz__zz_regVec_0 = regVec_1050;
      end
      12'b010000011011 : begin
        _zz__zz_regVec_0 = regVec_1051;
      end
      12'b010000011100 : begin
        _zz__zz_regVec_0 = regVec_1052;
      end
      12'b010000011101 : begin
        _zz__zz_regVec_0 = regVec_1053;
      end
      12'b010000011110 : begin
        _zz__zz_regVec_0 = regVec_1054;
      end
      12'b010000011111 : begin
        _zz__zz_regVec_0 = regVec_1055;
      end
      12'b010000100000 : begin
        _zz__zz_regVec_0 = regVec_1056;
      end
      12'b010000100001 : begin
        _zz__zz_regVec_0 = regVec_1057;
      end
      12'b010000100010 : begin
        _zz__zz_regVec_0 = regVec_1058;
      end
      12'b010000100011 : begin
        _zz__zz_regVec_0 = regVec_1059;
      end
      12'b010000100100 : begin
        _zz__zz_regVec_0 = regVec_1060;
      end
      12'b010000100101 : begin
        _zz__zz_regVec_0 = regVec_1061;
      end
      12'b010000100110 : begin
        _zz__zz_regVec_0 = regVec_1062;
      end
      12'b010000100111 : begin
        _zz__zz_regVec_0 = regVec_1063;
      end
      12'b010000101000 : begin
        _zz__zz_regVec_0 = regVec_1064;
      end
      12'b010000101001 : begin
        _zz__zz_regVec_0 = regVec_1065;
      end
      12'b010000101010 : begin
        _zz__zz_regVec_0 = regVec_1066;
      end
      12'b010000101011 : begin
        _zz__zz_regVec_0 = regVec_1067;
      end
      12'b010000101100 : begin
        _zz__zz_regVec_0 = regVec_1068;
      end
      12'b010000101101 : begin
        _zz__zz_regVec_0 = regVec_1069;
      end
      12'b010000101110 : begin
        _zz__zz_regVec_0 = regVec_1070;
      end
      12'b010000101111 : begin
        _zz__zz_regVec_0 = regVec_1071;
      end
      12'b010000110000 : begin
        _zz__zz_regVec_0 = regVec_1072;
      end
      12'b010000110001 : begin
        _zz__zz_regVec_0 = regVec_1073;
      end
      12'b010000110010 : begin
        _zz__zz_regVec_0 = regVec_1074;
      end
      12'b010000110011 : begin
        _zz__zz_regVec_0 = regVec_1075;
      end
      12'b010000110100 : begin
        _zz__zz_regVec_0 = regVec_1076;
      end
      12'b010000110101 : begin
        _zz__zz_regVec_0 = regVec_1077;
      end
      12'b010000110110 : begin
        _zz__zz_regVec_0 = regVec_1078;
      end
      12'b010000110111 : begin
        _zz__zz_regVec_0 = regVec_1079;
      end
      12'b010000111000 : begin
        _zz__zz_regVec_0 = regVec_1080;
      end
      12'b010000111001 : begin
        _zz__zz_regVec_0 = regVec_1081;
      end
      12'b010000111010 : begin
        _zz__zz_regVec_0 = regVec_1082;
      end
      12'b010000111011 : begin
        _zz__zz_regVec_0 = regVec_1083;
      end
      12'b010000111100 : begin
        _zz__zz_regVec_0 = regVec_1084;
      end
      12'b010000111101 : begin
        _zz__zz_regVec_0 = regVec_1085;
      end
      12'b010000111110 : begin
        _zz__zz_regVec_0 = regVec_1086;
      end
      12'b010000111111 : begin
        _zz__zz_regVec_0 = regVec_1087;
      end
      12'b010001000000 : begin
        _zz__zz_regVec_0 = regVec_1088;
      end
      12'b010001000001 : begin
        _zz__zz_regVec_0 = regVec_1089;
      end
      12'b010001000010 : begin
        _zz__zz_regVec_0 = regVec_1090;
      end
      12'b010001000011 : begin
        _zz__zz_regVec_0 = regVec_1091;
      end
      12'b010001000100 : begin
        _zz__zz_regVec_0 = regVec_1092;
      end
      12'b010001000101 : begin
        _zz__zz_regVec_0 = regVec_1093;
      end
      12'b010001000110 : begin
        _zz__zz_regVec_0 = regVec_1094;
      end
      12'b010001000111 : begin
        _zz__zz_regVec_0 = regVec_1095;
      end
      12'b010001001000 : begin
        _zz__zz_regVec_0 = regVec_1096;
      end
      12'b010001001001 : begin
        _zz__zz_regVec_0 = regVec_1097;
      end
      12'b010001001010 : begin
        _zz__zz_regVec_0 = regVec_1098;
      end
      12'b010001001011 : begin
        _zz__zz_regVec_0 = regVec_1099;
      end
      12'b010001001100 : begin
        _zz__zz_regVec_0 = regVec_1100;
      end
      12'b010001001101 : begin
        _zz__zz_regVec_0 = regVec_1101;
      end
      12'b010001001110 : begin
        _zz__zz_regVec_0 = regVec_1102;
      end
      12'b010001001111 : begin
        _zz__zz_regVec_0 = regVec_1103;
      end
      12'b010001010000 : begin
        _zz__zz_regVec_0 = regVec_1104;
      end
      12'b010001010001 : begin
        _zz__zz_regVec_0 = regVec_1105;
      end
      12'b010001010010 : begin
        _zz__zz_regVec_0 = regVec_1106;
      end
      12'b010001010011 : begin
        _zz__zz_regVec_0 = regVec_1107;
      end
      12'b010001010100 : begin
        _zz__zz_regVec_0 = regVec_1108;
      end
      12'b010001010101 : begin
        _zz__zz_regVec_0 = regVec_1109;
      end
      12'b010001010110 : begin
        _zz__zz_regVec_0 = regVec_1110;
      end
      12'b010001010111 : begin
        _zz__zz_regVec_0 = regVec_1111;
      end
      12'b010001011000 : begin
        _zz__zz_regVec_0 = regVec_1112;
      end
      12'b010001011001 : begin
        _zz__zz_regVec_0 = regVec_1113;
      end
      12'b010001011010 : begin
        _zz__zz_regVec_0 = regVec_1114;
      end
      12'b010001011011 : begin
        _zz__zz_regVec_0 = regVec_1115;
      end
      12'b010001011100 : begin
        _zz__zz_regVec_0 = regVec_1116;
      end
      12'b010001011101 : begin
        _zz__zz_regVec_0 = regVec_1117;
      end
      12'b010001011110 : begin
        _zz__zz_regVec_0 = regVec_1118;
      end
      12'b010001011111 : begin
        _zz__zz_regVec_0 = regVec_1119;
      end
      12'b010001100000 : begin
        _zz__zz_regVec_0 = regVec_1120;
      end
      12'b010001100001 : begin
        _zz__zz_regVec_0 = regVec_1121;
      end
      12'b010001100010 : begin
        _zz__zz_regVec_0 = regVec_1122;
      end
      12'b010001100011 : begin
        _zz__zz_regVec_0 = regVec_1123;
      end
      12'b010001100100 : begin
        _zz__zz_regVec_0 = regVec_1124;
      end
      12'b010001100101 : begin
        _zz__zz_regVec_0 = regVec_1125;
      end
      12'b010001100110 : begin
        _zz__zz_regVec_0 = regVec_1126;
      end
      12'b010001100111 : begin
        _zz__zz_regVec_0 = regVec_1127;
      end
      12'b010001101000 : begin
        _zz__zz_regVec_0 = regVec_1128;
      end
      12'b010001101001 : begin
        _zz__zz_regVec_0 = regVec_1129;
      end
      12'b010001101010 : begin
        _zz__zz_regVec_0 = regVec_1130;
      end
      12'b010001101011 : begin
        _zz__zz_regVec_0 = regVec_1131;
      end
      12'b010001101100 : begin
        _zz__zz_regVec_0 = regVec_1132;
      end
      12'b010001101101 : begin
        _zz__zz_regVec_0 = regVec_1133;
      end
      12'b010001101110 : begin
        _zz__zz_regVec_0 = regVec_1134;
      end
      12'b010001101111 : begin
        _zz__zz_regVec_0 = regVec_1135;
      end
      12'b010001110000 : begin
        _zz__zz_regVec_0 = regVec_1136;
      end
      12'b010001110001 : begin
        _zz__zz_regVec_0 = regVec_1137;
      end
      12'b010001110010 : begin
        _zz__zz_regVec_0 = regVec_1138;
      end
      12'b010001110011 : begin
        _zz__zz_regVec_0 = regVec_1139;
      end
      12'b010001110100 : begin
        _zz__zz_regVec_0 = regVec_1140;
      end
      12'b010001110101 : begin
        _zz__zz_regVec_0 = regVec_1141;
      end
      12'b010001110110 : begin
        _zz__zz_regVec_0 = regVec_1142;
      end
      12'b010001110111 : begin
        _zz__zz_regVec_0 = regVec_1143;
      end
      12'b010001111000 : begin
        _zz__zz_regVec_0 = regVec_1144;
      end
      12'b010001111001 : begin
        _zz__zz_regVec_0 = regVec_1145;
      end
      12'b010001111010 : begin
        _zz__zz_regVec_0 = regVec_1146;
      end
      12'b010001111011 : begin
        _zz__zz_regVec_0 = regVec_1147;
      end
      12'b010001111100 : begin
        _zz__zz_regVec_0 = regVec_1148;
      end
      12'b010001111101 : begin
        _zz__zz_regVec_0 = regVec_1149;
      end
      12'b010001111110 : begin
        _zz__zz_regVec_0 = regVec_1150;
      end
      12'b010001111111 : begin
        _zz__zz_regVec_0 = regVec_1151;
      end
      12'b010010000000 : begin
        _zz__zz_regVec_0 = regVec_1152;
      end
      12'b010010000001 : begin
        _zz__zz_regVec_0 = regVec_1153;
      end
      12'b010010000010 : begin
        _zz__zz_regVec_0 = regVec_1154;
      end
      12'b010010000011 : begin
        _zz__zz_regVec_0 = regVec_1155;
      end
      12'b010010000100 : begin
        _zz__zz_regVec_0 = regVec_1156;
      end
      12'b010010000101 : begin
        _zz__zz_regVec_0 = regVec_1157;
      end
      12'b010010000110 : begin
        _zz__zz_regVec_0 = regVec_1158;
      end
      12'b010010000111 : begin
        _zz__zz_regVec_0 = regVec_1159;
      end
      12'b010010001000 : begin
        _zz__zz_regVec_0 = regVec_1160;
      end
      12'b010010001001 : begin
        _zz__zz_regVec_0 = regVec_1161;
      end
      12'b010010001010 : begin
        _zz__zz_regVec_0 = regVec_1162;
      end
      12'b010010001011 : begin
        _zz__zz_regVec_0 = regVec_1163;
      end
      12'b010010001100 : begin
        _zz__zz_regVec_0 = regVec_1164;
      end
      12'b010010001101 : begin
        _zz__zz_regVec_0 = regVec_1165;
      end
      12'b010010001110 : begin
        _zz__zz_regVec_0 = regVec_1166;
      end
      12'b010010001111 : begin
        _zz__zz_regVec_0 = regVec_1167;
      end
      12'b010010010000 : begin
        _zz__zz_regVec_0 = regVec_1168;
      end
      12'b010010010001 : begin
        _zz__zz_regVec_0 = regVec_1169;
      end
      12'b010010010010 : begin
        _zz__zz_regVec_0 = regVec_1170;
      end
      12'b010010010011 : begin
        _zz__zz_regVec_0 = regVec_1171;
      end
      12'b010010010100 : begin
        _zz__zz_regVec_0 = regVec_1172;
      end
      12'b010010010101 : begin
        _zz__zz_regVec_0 = regVec_1173;
      end
      12'b010010010110 : begin
        _zz__zz_regVec_0 = regVec_1174;
      end
      12'b010010010111 : begin
        _zz__zz_regVec_0 = regVec_1175;
      end
      12'b010010011000 : begin
        _zz__zz_regVec_0 = regVec_1176;
      end
      12'b010010011001 : begin
        _zz__zz_regVec_0 = regVec_1177;
      end
      12'b010010011010 : begin
        _zz__zz_regVec_0 = regVec_1178;
      end
      12'b010010011011 : begin
        _zz__zz_regVec_0 = regVec_1179;
      end
      12'b010010011100 : begin
        _zz__zz_regVec_0 = regVec_1180;
      end
      12'b010010011101 : begin
        _zz__zz_regVec_0 = regVec_1181;
      end
      12'b010010011110 : begin
        _zz__zz_regVec_0 = regVec_1182;
      end
      12'b010010011111 : begin
        _zz__zz_regVec_0 = regVec_1183;
      end
      12'b010010100000 : begin
        _zz__zz_regVec_0 = regVec_1184;
      end
      12'b010010100001 : begin
        _zz__zz_regVec_0 = regVec_1185;
      end
      12'b010010100010 : begin
        _zz__zz_regVec_0 = regVec_1186;
      end
      12'b010010100011 : begin
        _zz__zz_regVec_0 = regVec_1187;
      end
      12'b010010100100 : begin
        _zz__zz_regVec_0 = regVec_1188;
      end
      12'b010010100101 : begin
        _zz__zz_regVec_0 = regVec_1189;
      end
      12'b010010100110 : begin
        _zz__zz_regVec_0 = regVec_1190;
      end
      12'b010010100111 : begin
        _zz__zz_regVec_0 = regVec_1191;
      end
      12'b010010101000 : begin
        _zz__zz_regVec_0 = regVec_1192;
      end
      12'b010010101001 : begin
        _zz__zz_regVec_0 = regVec_1193;
      end
      12'b010010101010 : begin
        _zz__zz_regVec_0 = regVec_1194;
      end
      12'b010010101011 : begin
        _zz__zz_regVec_0 = regVec_1195;
      end
      12'b010010101100 : begin
        _zz__zz_regVec_0 = regVec_1196;
      end
      12'b010010101101 : begin
        _zz__zz_regVec_0 = regVec_1197;
      end
      12'b010010101110 : begin
        _zz__zz_regVec_0 = regVec_1198;
      end
      12'b010010101111 : begin
        _zz__zz_regVec_0 = regVec_1199;
      end
      12'b010010110000 : begin
        _zz__zz_regVec_0 = regVec_1200;
      end
      12'b010010110001 : begin
        _zz__zz_regVec_0 = regVec_1201;
      end
      12'b010010110010 : begin
        _zz__zz_regVec_0 = regVec_1202;
      end
      12'b010010110011 : begin
        _zz__zz_regVec_0 = regVec_1203;
      end
      12'b010010110100 : begin
        _zz__zz_regVec_0 = regVec_1204;
      end
      12'b010010110101 : begin
        _zz__zz_regVec_0 = regVec_1205;
      end
      12'b010010110110 : begin
        _zz__zz_regVec_0 = regVec_1206;
      end
      12'b010010110111 : begin
        _zz__zz_regVec_0 = regVec_1207;
      end
      12'b010010111000 : begin
        _zz__zz_regVec_0 = regVec_1208;
      end
      12'b010010111001 : begin
        _zz__zz_regVec_0 = regVec_1209;
      end
      12'b010010111010 : begin
        _zz__zz_regVec_0 = regVec_1210;
      end
      12'b010010111011 : begin
        _zz__zz_regVec_0 = regVec_1211;
      end
      12'b010010111100 : begin
        _zz__zz_regVec_0 = regVec_1212;
      end
      12'b010010111101 : begin
        _zz__zz_regVec_0 = regVec_1213;
      end
      12'b010010111110 : begin
        _zz__zz_regVec_0 = regVec_1214;
      end
      12'b010010111111 : begin
        _zz__zz_regVec_0 = regVec_1215;
      end
      12'b010011000000 : begin
        _zz__zz_regVec_0 = regVec_1216;
      end
      12'b010011000001 : begin
        _zz__zz_regVec_0 = regVec_1217;
      end
      12'b010011000010 : begin
        _zz__zz_regVec_0 = regVec_1218;
      end
      12'b010011000011 : begin
        _zz__zz_regVec_0 = regVec_1219;
      end
      12'b010011000100 : begin
        _zz__zz_regVec_0 = regVec_1220;
      end
      12'b010011000101 : begin
        _zz__zz_regVec_0 = regVec_1221;
      end
      12'b010011000110 : begin
        _zz__zz_regVec_0 = regVec_1222;
      end
      12'b010011000111 : begin
        _zz__zz_regVec_0 = regVec_1223;
      end
      12'b010011001000 : begin
        _zz__zz_regVec_0 = regVec_1224;
      end
      12'b010011001001 : begin
        _zz__zz_regVec_0 = regVec_1225;
      end
      12'b010011001010 : begin
        _zz__zz_regVec_0 = regVec_1226;
      end
      12'b010011001011 : begin
        _zz__zz_regVec_0 = regVec_1227;
      end
      12'b010011001100 : begin
        _zz__zz_regVec_0 = regVec_1228;
      end
      12'b010011001101 : begin
        _zz__zz_regVec_0 = regVec_1229;
      end
      12'b010011001110 : begin
        _zz__zz_regVec_0 = regVec_1230;
      end
      12'b010011001111 : begin
        _zz__zz_regVec_0 = regVec_1231;
      end
      12'b010011010000 : begin
        _zz__zz_regVec_0 = regVec_1232;
      end
      12'b010011010001 : begin
        _zz__zz_regVec_0 = regVec_1233;
      end
      12'b010011010010 : begin
        _zz__zz_regVec_0 = regVec_1234;
      end
      12'b010011010011 : begin
        _zz__zz_regVec_0 = regVec_1235;
      end
      12'b010011010100 : begin
        _zz__zz_regVec_0 = regVec_1236;
      end
      12'b010011010101 : begin
        _zz__zz_regVec_0 = regVec_1237;
      end
      12'b010011010110 : begin
        _zz__zz_regVec_0 = regVec_1238;
      end
      12'b010011010111 : begin
        _zz__zz_regVec_0 = regVec_1239;
      end
      12'b010011011000 : begin
        _zz__zz_regVec_0 = regVec_1240;
      end
      12'b010011011001 : begin
        _zz__zz_regVec_0 = regVec_1241;
      end
      12'b010011011010 : begin
        _zz__zz_regVec_0 = regVec_1242;
      end
      12'b010011011011 : begin
        _zz__zz_regVec_0 = regVec_1243;
      end
      12'b010011011100 : begin
        _zz__zz_regVec_0 = regVec_1244;
      end
      12'b010011011101 : begin
        _zz__zz_regVec_0 = regVec_1245;
      end
      12'b010011011110 : begin
        _zz__zz_regVec_0 = regVec_1246;
      end
      12'b010011011111 : begin
        _zz__zz_regVec_0 = regVec_1247;
      end
      12'b010011100000 : begin
        _zz__zz_regVec_0 = regVec_1248;
      end
      12'b010011100001 : begin
        _zz__zz_regVec_0 = regVec_1249;
      end
      12'b010011100010 : begin
        _zz__zz_regVec_0 = regVec_1250;
      end
      12'b010011100011 : begin
        _zz__zz_regVec_0 = regVec_1251;
      end
      12'b010011100100 : begin
        _zz__zz_regVec_0 = regVec_1252;
      end
      12'b010011100101 : begin
        _zz__zz_regVec_0 = regVec_1253;
      end
      12'b010011100110 : begin
        _zz__zz_regVec_0 = regVec_1254;
      end
      12'b010011100111 : begin
        _zz__zz_regVec_0 = regVec_1255;
      end
      12'b010011101000 : begin
        _zz__zz_regVec_0 = regVec_1256;
      end
      12'b010011101001 : begin
        _zz__zz_regVec_0 = regVec_1257;
      end
      12'b010011101010 : begin
        _zz__zz_regVec_0 = regVec_1258;
      end
      12'b010011101011 : begin
        _zz__zz_regVec_0 = regVec_1259;
      end
      12'b010011101100 : begin
        _zz__zz_regVec_0 = regVec_1260;
      end
      12'b010011101101 : begin
        _zz__zz_regVec_0 = regVec_1261;
      end
      12'b010011101110 : begin
        _zz__zz_regVec_0 = regVec_1262;
      end
      12'b010011101111 : begin
        _zz__zz_regVec_0 = regVec_1263;
      end
      12'b010011110000 : begin
        _zz__zz_regVec_0 = regVec_1264;
      end
      12'b010011110001 : begin
        _zz__zz_regVec_0 = regVec_1265;
      end
      12'b010011110010 : begin
        _zz__zz_regVec_0 = regVec_1266;
      end
      12'b010011110011 : begin
        _zz__zz_regVec_0 = regVec_1267;
      end
      12'b010011110100 : begin
        _zz__zz_regVec_0 = regVec_1268;
      end
      12'b010011110101 : begin
        _zz__zz_regVec_0 = regVec_1269;
      end
      12'b010011110110 : begin
        _zz__zz_regVec_0 = regVec_1270;
      end
      12'b010011110111 : begin
        _zz__zz_regVec_0 = regVec_1271;
      end
      12'b010011111000 : begin
        _zz__zz_regVec_0 = regVec_1272;
      end
      12'b010011111001 : begin
        _zz__zz_regVec_0 = regVec_1273;
      end
      12'b010011111010 : begin
        _zz__zz_regVec_0 = regVec_1274;
      end
      12'b010011111011 : begin
        _zz__zz_regVec_0 = regVec_1275;
      end
      12'b010011111100 : begin
        _zz__zz_regVec_0 = regVec_1276;
      end
      12'b010011111101 : begin
        _zz__zz_regVec_0 = regVec_1277;
      end
      12'b010011111110 : begin
        _zz__zz_regVec_0 = regVec_1278;
      end
      12'b010011111111 : begin
        _zz__zz_regVec_0 = regVec_1279;
      end
      12'b010100000000 : begin
        _zz__zz_regVec_0 = regVec_1280;
      end
      12'b010100000001 : begin
        _zz__zz_regVec_0 = regVec_1281;
      end
      12'b010100000010 : begin
        _zz__zz_regVec_0 = regVec_1282;
      end
      12'b010100000011 : begin
        _zz__zz_regVec_0 = regVec_1283;
      end
      12'b010100000100 : begin
        _zz__zz_regVec_0 = regVec_1284;
      end
      12'b010100000101 : begin
        _zz__zz_regVec_0 = regVec_1285;
      end
      12'b010100000110 : begin
        _zz__zz_regVec_0 = regVec_1286;
      end
      12'b010100000111 : begin
        _zz__zz_regVec_0 = regVec_1287;
      end
      12'b010100001000 : begin
        _zz__zz_regVec_0 = regVec_1288;
      end
      12'b010100001001 : begin
        _zz__zz_regVec_0 = regVec_1289;
      end
      12'b010100001010 : begin
        _zz__zz_regVec_0 = regVec_1290;
      end
      12'b010100001011 : begin
        _zz__zz_regVec_0 = regVec_1291;
      end
      12'b010100001100 : begin
        _zz__zz_regVec_0 = regVec_1292;
      end
      12'b010100001101 : begin
        _zz__zz_regVec_0 = regVec_1293;
      end
      12'b010100001110 : begin
        _zz__zz_regVec_0 = regVec_1294;
      end
      12'b010100001111 : begin
        _zz__zz_regVec_0 = regVec_1295;
      end
      12'b010100010000 : begin
        _zz__zz_regVec_0 = regVec_1296;
      end
      12'b010100010001 : begin
        _zz__zz_regVec_0 = regVec_1297;
      end
      12'b010100010010 : begin
        _zz__zz_regVec_0 = regVec_1298;
      end
      12'b010100010011 : begin
        _zz__zz_regVec_0 = regVec_1299;
      end
      12'b010100010100 : begin
        _zz__zz_regVec_0 = regVec_1300;
      end
      12'b010100010101 : begin
        _zz__zz_regVec_0 = regVec_1301;
      end
      12'b010100010110 : begin
        _zz__zz_regVec_0 = regVec_1302;
      end
      12'b010100010111 : begin
        _zz__zz_regVec_0 = regVec_1303;
      end
      12'b010100011000 : begin
        _zz__zz_regVec_0 = regVec_1304;
      end
      12'b010100011001 : begin
        _zz__zz_regVec_0 = regVec_1305;
      end
      12'b010100011010 : begin
        _zz__zz_regVec_0 = regVec_1306;
      end
      12'b010100011011 : begin
        _zz__zz_regVec_0 = regVec_1307;
      end
      12'b010100011100 : begin
        _zz__zz_regVec_0 = regVec_1308;
      end
      12'b010100011101 : begin
        _zz__zz_regVec_0 = regVec_1309;
      end
      12'b010100011110 : begin
        _zz__zz_regVec_0 = regVec_1310;
      end
      12'b010100011111 : begin
        _zz__zz_regVec_0 = regVec_1311;
      end
      12'b010100100000 : begin
        _zz__zz_regVec_0 = regVec_1312;
      end
      12'b010100100001 : begin
        _zz__zz_regVec_0 = regVec_1313;
      end
      12'b010100100010 : begin
        _zz__zz_regVec_0 = regVec_1314;
      end
      12'b010100100011 : begin
        _zz__zz_regVec_0 = regVec_1315;
      end
      12'b010100100100 : begin
        _zz__zz_regVec_0 = regVec_1316;
      end
      12'b010100100101 : begin
        _zz__zz_regVec_0 = regVec_1317;
      end
      12'b010100100110 : begin
        _zz__zz_regVec_0 = regVec_1318;
      end
      12'b010100100111 : begin
        _zz__zz_regVec_0 = regVec_1319;
      end
      12'b010100101000 : begin
        _zz__zz_regVec_0 = regVec_1320;
      end
      12'b010100101001 : begin
        _zz__zz_regVec_0 = regVec_1321;
      end
      12'b010100101010 : begin
        _zz__zz_regVec_0 = regVec_1322;
      end
      12'b010100101011 : begin
        _zz__zz_regVec_0 = regVec_1323;
      end
      12'b010100101100 : begin
        _zz__zz_regVec_0 = regVec_1324;
      end
      12'b010100101101 : begin
        _zz__zz_regVec_0 = regVec_1325;
      end
      12'b010100101110 : begin
        _zz__zz_regVec_0 = regVec_1326;
      end
      12'b010100101111 : begin
        _zz__zz_regVec_0 = regVec_1327;
      end
      12'b010100110000 : begin
        _zz__zz_regVec_0 = regVec_1328;
      end
      12'b010100110001 : begin
        _zz__zz_regVec_0 = regVec_1329;
      end
      12'b010100110010 : begin
        _zz__zz_regVec_0 = regVec_1330;
      end
      12'b010100110011 : begin
        _zz__zz_regVec_0 = regVec_1331;
      end
      12'b010100110100 : begin
        _zz__zz_regVec_0 = regVec_1332;
      end
      12'b010100110101 : begin
        _zz__zz_regVec_0 = regVec_1333;
      end
      12'b010100110110 : begin
        _zz__zz_regVec_0 = regVec_1334;
      end
      12'b010100110111 : begin
        _zz__zz_regVec_0 = regVec_1335;
      end
      12'b010100111000 : begin
        _zz__zz_regVec_0 = regVec_1336;
      end
      12'b010100111001 : begin
        _zz__zz_regVec_0 = regVec_1337;
      end
      12'b010100111010 : begin
        _zz__zz_regVec_0 = regVec_1338;
      end
      12'b010100111011 : begin
        _zz__zz_regVec_0 = regVec_1339;
      end
      12'b010100111100 : begin
        _zz__zz_regVec_0 = regVec_1340;
      end
      12'b010100111101 : begin
        _zz__zz_regVec_0 = regVec_1341;
      end
      12'b010100111110 : begin
        _zz__zz_regVec_0 = regVec_1342;
      end
      12'b010100111111 : begin
        _zz__zz_regVec_0 = regVec_1343;
      end
      12'b010101000000 : begin
        _zz__zz_regVec_0 = regVec_1344;
      end
      12'b010101000001 : begin
        _zz__zz_regVec_0 = regVec_1345;
      end
      12'b010101000010 : begin
        _zz__zz_regVec_0 = regVec_1346;
      end
      12'b010101000011 : begin
        _zz__zz_regVec_0 = regVec_1347;
      end
      12'b010101000100 : begin
        _zz__zz_regVec_0 = regVec_1348;
      end
      12'b010101000101 : begin
        _zz__zz_regVec_0 = regVec_1349;
      end
      12'b010101000110 : begin
        _zz__zz_regVec_0 = regVec_1350;
      end
      12'b010101000111 : begin
        _zz__zz_regVec_0 = regVec_1351;
      end
      12'b010101001000 : begin
        _zz__zz_regVec_0 = regVec_1352;
      end
      12'b010101001001 : begin
        _zz__zz_regVec_0 = regVec_1353;
      end
      12'b010101001010 : begin
        _zz__zz_regVec_0 = regVec_1354;
      end
      12'b010101001011 : begin
        _zz__zz_regVec_0 = regVec_1355;
      end
      12'b010101001100 : begin
        _zz__zz_regVec_0 = regVec_1356;
      end
      12'b010101001101 : begin
        _zz__zz_regVec_0 = regVec_1357;
      end
      12'b010101001110 : begin
        _zz__zz_regVec_0 = regVec_1358;
      end
      12'b010101001111 : begin
        _zz__zz_regVec_0 = regVec_1359;
      end
      12'b010101010000 : begin
        _zz__zz_regVec_0 = regVec_1360;
      end
      12'b010101010001 : begin
        _zz__zz_regVec_0 = regVec_1361;
      end
      12'b010101010010 : begin
        _zz__zz_regVec_0 = regVec_1362;
      end
      12'b010101010011 : begin
        _zz__zz_regVec_0 = regVec_1363;
      end
      12'b010101010100 : begin
        _zz__zz_regVec_0 = regVec_1364;
      end
      12'b010101010101 : begin
        _zz__zz_regVec_0 = regVec_1365;
      end
      12'b010101010110 : begin
        _zz__zz_regVec_0 = regVec_1366;
      end
      12'b010101010111 : begin
        _zz__zz_regVec_0 = regVec_1367;
      end
      12'b010101011000 : begin
        _zz__zz_regVec_0 = regVec_1368;
      end
      12'b010101011001 : begin
        _zz__zz_regVec_0 = regVec_1369;
      end
      12'b010101011010 : begin
        _zz__zz_regVec_0 = regVec_1370;
      end
      12'b010101011011 : begin
        _zz__zz_regVec_0 = regVec_1371;
      end
      12'b010101011100 : begin
        _zz__zz_regVec_0 = regVec_1372;
      end
      12'b010101011101 : begin
        _zz__zz_regVec_0 = regVec_1373;
      end
      12'b010101011110 : begin
        _zz__zz_regVec_0 = regVec_1374;
      end
      12'b010101011111 : begin
        _zz__zz_regVec_0 = regVec_1375;
      end
      12'b010101100000 : begin
        _zz__zz_regVec_0 = regVec_1376;
      end
      12'b010101100001 : begin
        _zz__zz_regVec_0 = regVec_1377;
      end
      12'b010101100010 : begin
        _zz__zz_regVec_0 = regVec_1378;
      end
      12'b010101100011 : begin
        _zz__zz_regVec_0 = regVec_1379;
      end
      12'b010101100100 : begin
        _zz__zz_regVec_0 = regVec_1380;
      end
      12'b010101100101 : begin
        _zz__zz_regVec_0 = regVec_1381;
      end
      12'b010101100110 : begin
        _zz__zz_regVec_0 = regVec_1382;
      end
      12'b010101100111 : begin
        _zz__zz_regVec_0 = regVec_1383;
      end
      12'b010101101000 : begin
        _zz__zz_regVec_0 = regVec_1384;
      end
      12'b010101101001 : begin
        _zz__zz_regVec_0 = regVec_1385;
      end
      12'b010101101010 : begin
        _zz__zz_regVec_0 = regVec_1386;
      end
      12'b010101101011 : begin
        _zz__zz_regVec_0 = regVec_1387;
      end
      12'b010101101100 : begin
        _zz__zz_regVec_0 = regVec_1388;
      end
      12'b010101101101 : begin
        _zz__zz_regVec_0 = regVec_1389;
      end
      12'b010101101110 : begin
        _zz__zz_regVec_0 = regVec_1390;
      end
      12'b010101101111 : begin
        _zz__zz_regVec_0 = regVec_1391;
      end
      12'b010101110000 : begin
        _zz__zz_regVec_0 = regVec_1392;
      end
      12'b010101110001 : begin
        _zz__zz_regVec_0 = regVec_1393;
      end
      12'b010101110010 : begin
        _zz__zz_regVec_0 = regVec_1394;
      end
      12'b010101110011 : begin
        _zz__zz_regVec_0 = regVec_1395;
      end
      12'b010101110100 : begin
        _zz__zz_regVec_0 = regVec_1396;
      end
      12'b010101110101 : begin
        _zz__zz_regVec_0 = regVec_1397;
      end
      12'b010101110110 : begin
        _zz__zz_regVec_0 = regVec_1398;
      end
      12'b010101110111 : begin
        _zz__zz_regVec_0 = regVec_1399;
      end
      12'b010101111000 : begin
        _zz__zz_regVec_0 = regVec_1400;
      end
      12'b010101111001 : begin
        _zz__zz_regVec_0 = regVec_1401;
      end
      12'b010101111010 : begin
        _zz__zz_regVec_0 = regVec_1402;
      end
      12'b010101111011 : begin
        _zz__zz_regVec_0 = regVec_1403;
      end
      12'b010101111100 : begin
        _zz__zz_regVec_0 = regVec_1404;
      end
      12'b010101111101 : begin
        _zz__zz_regVec_0 = regVec_1405;
      end
      12'b010101111110 : begin
        _zz__zz_regVec_0 = regVec_1406;
      end
      12'b010101111111 : begin
        _zz__zz_regVec_0 = regVec_1407;
      end
      12'b010110000000 : begin
        _zz__zz_regVec_0 = regVec_1408;
      end
      12'b010110000001 : begin
        _zz__zz_regVec_0 = regVec_1409;
      end
      12'b010110000010 : begin
        _zz__zz_regVec_0 = regVec_1410;
      end
      12'b010110000011 : begin
        _zz__zz_regVec_0 = regVec_1411;
      end
      12'b010110000100 : begin
        _zz__zz_regVec_0 = regVec_1412;
      end
      12'b010110000101 : begin
        _zz__zz_regVec_0 = regVec_1413;
      end
      12'b010110000110 : begin
        _zz__zz_regVec_0 = regVec_1414;
      end
      12'b010110000111 : begin
        _zz__zz_regVec_0 = regVec_1415;
      end
      12'b010110001000 : begin
        _zz__zz_regVec_0 = regVec_1416;
      end
      12'b010110001001 : begin
        _zz__zz_regVec_0 = regVec_1417;
      end
      12'b010110001010 : begin
        _zz__zz_regVec_0 = regVec_1418;
      end
      12'b010110001011 : begin
        _zz__zz_regVec_0 = regVec_1419;
      end
      12'b010110001100 : begin
        _zz__zz_regVec_0 = regVec_1420;
      end
      12'b010110001101 : begin
        _zz__zz_regVec_0 = regVec_1421;
      end
      12'b010110001110 : begin
        _zz__zz_regVec_0 = regVec_1422;
      end
      12'b010110001111 : begin
        _zz__zz_regVec_0 = regVec_1423;
      end
      12'b010110010000 : begin
        _zz__zz_regVec_0 = regVec_1424;
      end
      12'b010110010001 : begin
        _zz__zz_regVec_0 = regVec_1425;
      end
      12'b010110010010 : begin
        _zz__zz_regVec_0 = regVec_1426;
      end
      12'b010110010011 : begin
        _zz__zz_regVec_0 = regVec_1427;
      end
      12'b010110010100 : begin
        _zz__zz_regVec_0 = regVec_1428;
      end
      12'b010110010101 : begin
        _zz__zz_regVec_0 = regVec_1429;
      end
      12'b010110010110 : begin
        _zz__zz_regVec_0 = regVec_1430;
      end
      12'b010110010111 : begin
        _zz__zz_regVec_0 = regVec_1431;
      end
      12'b010110011000 : begin
        _zz__zz_regVec_0 = regVec_1432;
      end
      12'b010110011001 : begin
        _zz__zz_regVec_0 = regVec_1433;
      end
      12'b010110011010 : begin
        _zz__zz_regVec_0 = regVec_1434;
      end
      12'b010110011011 : begin
        _zz__zz_regVec_0 = regVec_1435;
      end
      12'b010110011100 : begin
        _zz__zz_regVec_0 = regVec_1436;
      end
      12'b010110011101 : begin
        _zz__zz_regVec_0 = regVec_1437;
      end
      12'b010110011110 : begin
        _zz__zz_regVec_0 = regVec_1438;
      end
      12'b010110011111 : begin
        _zz__zz_regVec_0 = regVec_1439;
      end
      12'b010110100000 : begin
        _zz__zz_regVec_0 = regVec_1440;
      end
      12'b010110100001 : begin
        _zz__zz_regVec_0 = regVec_1441;
      end
      12'b010110100010 : begin
        _zz__zz_regVec_0 = regVec_1442;
      end
      12'b010110100011 : begin
        _zz__zz_regVec_0 = regVec_1443;
      end
      12'b010110100100 : begin
        _zz__zz_regVec_0 = regVec_1444;
      end
      12'b010110100101 : begin
        _zz__zz_regVec_0 = regVec_1445;
      end
      12'b010110100110 : begin
        _zz__zz_regVec_0 = regVec_1446;
      end
      12'b010110100111 : begin
        _zz__zz_regVec_0 = regVec_1447;
      end
      12'b010110101000 : begin
        _zz__zz_regVec_0 = regVec_1448;
      end
      12'b010110101001 : begin
        _zz__zz_regVec_0 = regVec_1449;
      end
      12'b010110101010 : begin
        _zz__zz_regVec_0 = regVec_1450;
      end
      12'b010110101011 : begin
        _zz__zz_regVec_0 = regVec_1451;
      end
      12'b010110101100 : begin
        _zz__zz_regVec_0 = regVec_1452;
      end
      12'b010110101101 : begin
        _zz__zz_regVec_0 = regVec_1453;
      end
      12'b010110101110 : begin
        _zz__zz_regVec_0 = regVec_1454;
      end
      12'b010110101111 : begin
        _zz__zz_regVec_0 = regVec_1455;
      end
      12'b010110110000 : begin
        _zz__zz_regVec_0 = regVec_1456;
      end
      12'b010110110001 : begin
        _zz__zz_regVec_0 = regVec_1457;
      end
      12'b010110110010 : begin
        _zz__zz_regVec_0 = regVec_1458;
      end
      12'b010110110011 : begin
        _zz__zz_regVec_0 = regVec_1459;
      end
      12'b010110110100 : begin
        _zz__zz_regVec_0 = regVec_1460;
      end
      12'b010110110101 : begin
        _zz__zz_regVec_0 = regVec_1461;
      end
      12'b010110110110 : begin
        _zz__zz_regVec_0 = regVec_1462;
      end
      12'b010110110111 : begin
        _zz__zz_regVec_0 = regVec_1463;
      end
      12'b010110111000 : begin
        _zz__zz_regVec_0 = regVec_1464;
      end
      12'b010110111001 : begin
        _zz__zz_regVec_0 = regVec_1465;
      end
      12'b010110111010 : begin
        _zz__zz_regVec_0 = regVec_1466;
      end
      12'b010110111011 : begin
        _zz__zz_regVec_0 = regVec_1467;
      end
      12'b010110111100 : begin
        _zz__zz_regVec_0 = regVec_1468;
      end
      12'b010110111101 : begin
        _zz__zz_regVec_0 = regVec_1469;
      end
      12'b010110111110 : begin
        _zz__zz_regVec_0 = regVec_1470;
      end
      12'b010110111111 : begin
        _zz__zz_regVec_0 = regVec_1471;
      end
      12'b010111000000 : begin
        _zz__zz_regVec_0 = regVec_1472;
      end
      12'b010111000001 : begin
        _zz__zz_regVec_0 = regVec_1473;
      end
      12'b010111000010 : begin
        _zz__zz_regVec_0 = regVec_1474;
      end
      12'b010111000011 : begin
        _zz__zz_regVec_0 = regVec_1475;
      end
      12'b010111000100 : begin
        _zz__zz_regVec_0 = regVec_1476;
      end
      12'b010111000101 : begin
        _zz__zz_regVec_0 = regVec_1477;
      end
      12'b010111000110 : begin
        _zz__zz_regVec_0 = regVec_1478;
      end
      12'b010111000111 : begin
        _zz__zz_regVec_0 = regVec_1479;
      end
      12'b010111001000 : begin
        _zz__zz_regVec_0 = regVec_1480;
      end
      12'b010111001001 : begin
        _zz__zz_regVec_0 = regVec_1481;
      end
      12'b010111001010 : begin
        _zz__zz_regVec_0 = regVec_1482;
      end
      12'b010111001011 : begin
        _zz__zz_regVec_0 = regVec_1483;
      end
      12'b010111001100 : begin
        _zz__zz_regVec_0 = regVec_1484;
      end
      12'b010111001101 : begin
        _zz__zz_regVec_0 = regVec_1485;
      end
      12'b010111001110 : begin
        _zz__zz_regVec_0 = regVec_1486;
      end
      12'b010111001111 : begin
        _zz__zz_regVec_0 = regVec_1487;
      end
      12'b010111010000 : begin
        _zz__zz_regVec_0 = regVec_1488;
      end
      12'b010111010001 : begin
        _zz__zz_regVec_0 = regVec_1489;
      end
      12'b010111010010 : begin
        _zz__zz_regVec_0 = regVec_1490;
      end
      12'b010111010011 : begin
        _zz__zz_regVec_0 = regVec_1491;
      end
      12'b010111010100 : begin
        _zz__zz_regVec_0 = regVec_1492;
      end
      12'b010111010101 : begin
        _zz__zz_regVec_0 = regVec_1493;
      end
      12'b010111010110 : begin
        _zz__zz_regVec_0 = regVec_1494;
      end
      12'b010111010111 : begin
        _zz__zz_regVec_0 = regVec_1495;
      end
      12'b010111011000 : begin
        _zz__zz_regVec_0 = regVec_1496;
      end
      12'b010111011001 : begin
        _zz__zz_regVec_0 = regVec_1497;
      end
      12'b010111011010 : begin
        _zz__zz_regVec_0 = regVec_1498;
      end
      12'b010111011011 : begin
        _zz__zz_regVec_0 = regVec_1499;
      end
      12'b010111011100 : begin
        _zz__zz_regVec_0 = regVec_1500;
      end
      12'b010111011101 : begin
        _zz__zz_regVec_0 = regVec_1501;
      end
      12'b010111011110 : begin
        _zz__zz_regVec_0 = regVec_1502;
      end
      12'b010111011111 : begin
        _zz__zz_regVec_0 = regVec_1503;
      end
      12'b010111100000 : begin
        _zz__zz_regVec_0 = regVec_1504;
      end
      12'b010111100001 : begin
        _zz__zz_regVec_0 = regVec_1505;
      end
      12'b010111100010 : begin
        _zz__zz_regVec_0 = regVec_1506;
      end
      12'b010111100011 : begin
        _zz__zz_regVec_0 = regVec_1507;
      end
      12'b010111100100 : begin
        _zz__zz_regVec_0 = regVec_1508;
      end
      12'b010111100101 : begin
        _zz__zz_regVec_0 = regVec_1509;
      end
      12'b010111100110 : begin
        _zz__zz_regVec_0 = regVec_1510;
      end
      12'b010111100111 : begin
        _zz__zz_regVec_0 = regVec_1511;
      end
      12'b010111101000 : begin
        _zz__zz_regVec_0 = regVec_1512;
      end
      12'b010111101001 : begin
        _zz__zz_regVec_0 = regVec_1513;
      end
      12'b010111101010 : begin
        _zz__zz_regVec_0 = regVec_1514;
      end
      12'b010111101011 : begin
        _zz__zz_regVec_0 = regVec_1515;
      end
      12'b010111101100 : begin
        _zz__zz_regVec_0 = regVec_1516;
      end
      12'b010111101101 : begin
        _zz__zz_regVec_0 = regVec_1517;
      end
      12'b010111101110 : begin
        _zz__zz_regVec_0 = regVec_1518;
      end
      12'b010111101111 : begin
        _zz__zz_regVec_0 = regVec_1519;
      end
      12'b010111110000 : begin
        _zz__zz_regVec_0 = regVec_1520;
      end
      12'b010111110001 : begin
        _zz__zz_regVec_0 = regVec_1521;
      end
      12'b010111110010 : begin
        _zz__zz_regVec_0 = regVec_1522;
      end
      12'b010111110011 : begin
        _zz__zz_regVec_0 = regVec_1523;
      end
      12'b010111110100 : begin
        _zz__zz_regVec_0 = regVec_1524;
      end
      12'b010111110101 : begin
        _zz__zz_regVec_0 = regVec_1525;
      end
      12'b010111110110 : begin
        _zz__zz_regVec_0 = regVec_1526;
      end
      12'b010111110111 : begin
        _zz__zz_regVec_0 = regVec_1527;
      end
      12'b010111111000 : begin
        _zz__zz_regVec_0 = regVec_1528;
      end
      12'b010111111001 : begin
        _zz__zz_regVec_0 = regVec_1529;
      end
      12'b010111111010 : begin
        _zz__zz_regVec_0 = regVec_1530;
      end
      12'b010111111011 : begin
        _zz__zz_regVec_0 = regVec_1531;
      end
      12'b010111111100 : begin
        _zz__zz_regVec_0 = regVec_1532;
      end
      12'b010111111101 : begin
        _zz__zz_regVec_0 = regVec_1533;
      end
      12'b010111111110 : begin
        _zz__zz_regVec_0 = regVec_1534;
      end
      12'b010111111111 : begin
        _zz__zz_regVec_0 = regVec_1535;
      end
      12'b011000000000 : begin
        _zz__zz_regVec_0 = regVec_1536;
      end
      12'b011000000001 : begin
        _zz__zz_regVec_0 = regVec_1537;
      end
      12'b011000000010 : begin
        _zz__zz_regVec_0 = regVec_1538;
      end
      12'b011000000011 : begin
        _zz__zz_regVec_0 = regVec_1539;
      end
      12'b011000000100 : begin
        _zz__zz_regVec_0 = regVec_1540;
      end
      12'b011000000101 : begin
        _zz__zz_regVec_0 = regVec_1541;
      end
      12'b011000000110 : begin
        _zz__zz_regVec_0 = regVec_1542;
      end
      12'b011000000111 : begin
        _zz__zz_regVec_0 = regVec_1543;
      end
      12'b011000001000 : begin
        _zz__zz_regVec_0 = regVec_1544;
      end
      12'b011000001001 : begin
        _zz__zz_regVec_0 = regVec_1545;
      end
      12'b011000001010 : begin
        _zz__zz_regVec_0 = regVec_1546;
      end
      12'b011000001011 : begin
        _zz__zz_regVec_0 = regVec_1547;
      end
      12'b011000001100 : begin
        _zz__zz_regVec_0 = regVec_1548;
      end
      12'b011000001101 : begin
        _zz__zz_regVec_0 = regVec_1549;
      end
      12'b011000001110 : begin
        _zz__zz_regVec_0 = regVec_1550;
      end
      12'b011000001111 : begin
        _zz__zz_regVec_0 = regVec_1551;
      end
      12'b011000010000 : begin
        _zz__zz_regVec_0 = regVec_1552;
      end
      12'b011000010001 : begin
        _zz__zz_regVec_0 = regVec_1553;
      end
      12'b011000010010 : begin
        _zz__zz_regVec_0 = regVec_1554;
      end
      12'b011000010011 : begin
        _zz__zz_regVec_0 = regVec_1555;
      end
      12'b011000010100 : begin
        _zz__zz_regVec_0 = regVec_1556;
      end
      12'b011000010101 : begin
        _zz__zz_regVec_0 = regVec_1557;
      end
      12'b011000010110 : begin
        _zz__zz_regVec_0 = regVec_1558;
      end
      12'b011000010111 : begin
        _zz__zz_regVec_0 = regVec_1559;
      end
      12'b011000011000 : begin
        _zz__zz_regVec_0 = regVec_1560;
      end
      12'b011000011001 : begin
        _zz__zz_regVec_0 = regVec_1561;
      end
      12'b011000011010 : begin
        _zz__zz_regVec_0 = regVec_1562;
      end
      12'b011000011011 : begin
        _zz__zz_regVec_0 = regVec_1563;
      end
      12'b011000011100 : begin
        _zz__zz_regVec_0 = regVec_1564;
      end
      12'b011000011101 : begin
        _zz__zz_regVec_0 = regVec_1565;
      end
      12'b011000011110 : begin
        _zz__zz_regVec_0 = regVec_1566;
      end
      12'b011000011111 : begin
        _zz__zz_regVec_0 = regVec_1567;
      end
      12'b011000100000 : begin
        _zz__zz_regVec_0 = regVec_1568;
      end
      12'b011000100001 : begin
        _zz__zz_regVec_0 = regVec_1569;
      end
      12'b011000100010 : begin
        _zz__zz_regVec_0 = regVec_1570;
      end
      12'b011000100011 : begin
        _zz__zz_regVec_0 = regVec_1571;
      end
      12'b011000100100 : begin
        _zz__zz_regVec_0 = regVec_1572;
      end
      12'b011000100101 : begin
        _zz__zz_regVec_0 = regVec_1573;
      end
      12'b011000100110 : begin
        _zz__zz_regVec_0 = regVec_1574;
      end
      12'b011000100111 : begin
        _zz__zz_regVec_0 = regVec_1575;
      end
      12'b011000101000 : begin
        _zz__zz_regVec_0 = regVec_1576;
      end
      12'b011000101001 : begin
        _zz__zz_regVec_0 = regVec_1577;
      end
      12'b011000101010 : begin
        _zz__zz_regVec_0 = regVec_1578;
      end
      12'b011000101011 : begin
        _zz__zz_regVec_0 = regVec_1579;
      end
      12'b011000101100 : begin
        _zz__zz_regVec_0 = regVec_1580;
      end
      12'b011000101101 : begin
        _zz__zz_regVec_0 = regVec_1581;
      end
      12'b011000101110 : begin
        _zz__zz_regVec_0 = regVec_1582;
      end
      12'b011000101111 : begin
        _zz__zz_regVec_0 = regVec_1583;
      end
      12'b011000110000 : begin
        _zz__zz_regVec_0 = regVec_1584;
      end
      12'b011000110001 : begin
        _zz__zz_regVec_0 = regVec_1585;
      end
      12'b011000110010 : begin
        _zz__zz_regVec_0 = regVec_1586;
      end
      12'b011000110011 : begin
        _zz__zz_regVec_0 = regVec_1587;
      end
      12'b011000110100 : begin
        _zz__zz_regVec_0 = regVec_1588;
      end
      12'b011000110101 : begin
        _zz__zz_regVec_0 = regVec_1589;
      end
      12'b011000110110 : begin
        _zz__zz_regVec_0 = regVec_1590;
      end
      12'b011000110111 : begin
        _zz__zz_regVec_0 = regVec_1591;
      end
      12'b011000111000 : begin
        _zz__zz_regVec_0 = regVec_1592;
      end
      12'b011000111001 : begin
        _zz__zz_regVec_0 = regVec_1593;
      end
      12'b011000111010 : begin
        _zz__zz_regVec_0 = regVec_1594;
      end
      12'b011000111011 : begin
        _zz__zz_regVec_0 = regVec_1595;
      end
      12'b011000111100 : begin
        _zz__zz_regVec_0 = regVec_1596;
      end
      12'b011000111101 : begin
        _zz__zz_regVec_0 = regVec_1597;
      end
      12'b011000111110 : begin
        _zz__zz_regVec_0 = regVec_1598;
      end
      12'b011000111111 : begin
        _zz__zz_regVec_0 = regVec_1599;
      end
      12'b011001000000 : begin
        _zz__zz_regVec_0 = regVec_1600;
      end
      12'b011001000001 : begin
        _zz__zz_regVec_0 = regVec_1601;
      end
      12'b011001000010 : begin
        _zz__zz_regVec_0 = regVec_1602;
      end
      12'b011001000011 : begin
        _zz__zz_regVec_0 = regVec_1603;
      end
      12'b011001000100 : begin
        _zz__zz_regVec_0 = regVec_1604;
      end
      12'b011001000101 : begin
        _zz__zz_regVec_0 = regVec_1605;
      end
      12'b011001000110 : begin
        _zz__zz_regVec_0 = regVec_1606;
      end
      12'b011001000111 : begin
        _zz__zz_regVec_0 = regVec_1607;
      end
      12'b011001001000 : begin
        _zz__zz_regVec_0 = regVec_1608;
      end
      12'b011001001001 : begin
        _zz__zz_regVec_0 = regVec_1609;
      end
      12'b011001001010 : begin
        _zz__zz_regVec_0 = regVec_1610;
      end
      12'b011001001011 : begin
        _zz__zz_regVec_0 = regVec_1611;
      end
      12'b011001001100 : begin
        _zz__zz_regVec_0 = regVec_1612;
      end
      12'b011001001101 : begin
        _zz__zz_regVec_0 = regVec_1613;
      end
      12'b011001001110 : begin
        _zz__zz_regVec_0 = regVec_1614;
      end
      12'b011001001111 : begin
        _zz__zz_regVec_0 = regVec_1615;
      end
      12'b011001010000 : begin
        _zz__zz_regVec_0 = regVec_1616;
      end
      12'b011001010001 : begin
        _zz__zz_regVec_0 = regVec_1617;
      end
      12'b011001010010 : begin
        _zz__zz_regVec_0 = regVec_1618;
      end
      12'b011001010011 : begin
        _zz__zz_regVec_0 = regVec_1619;
      end
      12'b011001010100 : begin
        _zz__zz_regVec_0 = regVec_1620;
      end
      12'b011001010101 : begin
        _zz__zz_regVec_0 = regVec_1621;
      end
      12'b011001010110 : begin
        _zz__zz_regVec_0 = regVec_1622;
      end
      12'b011001010111 : begin
        _zz__zz_regVec_0 = regVec_1623;
      end
      12'b011001011000 : begin
        _zz__zz_regVec_0 = regVec_1624;
      end
      12'b011001011001 : begin
        _zz__zz_regVec_0 = regVec_1625;
      end
      12'b011001011010 : begin
        _zz__zz_regVec_0 = regVec_1626;
      end
      12'b011001011011 : begin
        _zz__zz_regVec_0 = regVec_1627;
      end
      12'b011001011100 : begin
        _zz__zz_regVec_0 = regVec_1628;
      end
      12'b011001011101 : begin
        _zz__zz_regVec_0 = regVec_1629;
      end
      12'b011001011110 : begin
        _zz__zz_regVec_0 = regVec_1630;
      end
      12'b011001011111 : begin
        _zz__zz_regVec_0 = regVec_1631;
      end
      12'b011001100000 : begin
        _zz__zz_regVec_0 = regVec_1632;
      end
      12'b011001100001 : begin
        _zz__zz_regVec_0 = regVec_1633;
      end
      12'b011001100010 : begin
        _zz__zz_regVec_0 = regVec_1634;
      end
      12'b011001100011 : begin
        _zz__zz_regVec_0 = regVec_1635;
      end
      12'b011001100100 : begin
        _zz__zz_regVec_0 = regVec_1636;
      end
      12'b011001100101 : begin
        _zz__zz_regVec_0 = regVec_1637;
      end
      12'b011001100110 : begin
        _zz__zz_regVec_0 = regVec_1638;
      end
      12'b011001100111 : begin
        _zz__zz_regVec_0 = regVec_1639;
      end
      12'b011001101000 : begin
        _zz__zz_regVec_0 = regVec_1640;
      end
      12'b011001101001 : begin
        _zz__zz_regVec_0 = regVec_1641;
      end
      12'b011001101010 : begin
        _zz__zz_regVec_0 = regVec_1642;
      end
      12'b011001101011 : begin
        _zz__zz_regVec_0 = regVec_1643;
      end
      12'b011001101100 : begin
        _zz__zz_regVec_0 = regVec_1644;
      end
      12'b011001101101 : begin
        _zz__zz_regVec_0 = regVec_1645;
      end
      12'b011001101110 : begin
        _zz__zz_regVec_0 = regVec_1646;
      end
      12'b011001101111 : begin
        _zz__zz_regVec_0 = regVec_1647;
      end
      12'b011001110000 : begin
        _zz__zz_regVec_0 = regVec_1648;
      end
      12'b011001110001 : begin
        _zz__zz_regVec_0 = regVec_1649;
      end
      12'b011001110010 : begin
        _zz__zz_regVec_0 = regVec_1650;
      end
      12'b011001110011 : begin
        _zz__zz_regVec_0 = regVec_1651;
      end
      12'b011001110100 : begin
        _zz__zz_regVec_0 = regVec_1652;
      end
      12'b011001110101 : begin
        _zz__zz_regVec_0 = regVec_1653;
      end
      12'b011001110110 : begin
        _zz__zz_regVec_0 = regVec_1654;
      end
      12'b011001110111 : begin
        _zz__zz_regVec_0 = regVec_1655;
      end
      12'b011001111000 : begin
        _zz__zz_regVec_0 = regVec_1656;
      end
      12'b011001111001 : begin
        _zz__zz_regVec_0 = regVec_1657;
      end
      12'b011001111010 : begin
        _zz__zz_regVec_0 = regVec_1658;
      end
      12'b011001111011 : begin
        _zz__zz_regVec_0 = regVec_1659;
      end
      12'b011001111100 : begin
        _zz__zz_regVec_0 = regVec_1660;
      end
      12'b011001111101 : begin
        _zz__zz_regVec_0 = regVec_1661;
      end
      12'b011001111110 : begin
        _zz__zz_regVec_0 = regVec_1662;
      end
      12'b011001111111 : begin
        _zz__zz_regVec_0 = regVec_1663;
      end
      12'b011010000000 : begin
        _zz__zz_regVec_0 = regVec_1664;
      end
      12'b011010000001 : begin
        _zz__zz_regVec_0 = regVec_1665;
      end
      12'b011010000010 : begin
        _zz__zz_regVec_0 = regVec_1666;
      end
      12'b011010000011 : begin
        _zz__zz_regVec_0 = regVec_1667;
      end
      12'b011010000100 : begin
        _zz__zz_regVec_0 = regVec_1668;
      end
      12'b011010000101 : begin
        _zz__zz_regVec_0 = regVec_1669;
      end
      12'b011010000110 : begin
        _zz__zz_regVec_0 = regVec_1670;
      end
      12'b011010000111 : begin
        _zz__zz_regVec_0 = regVec_1671;
      end
      12'b011010001000 : begin
        _zz__zz_regVec_0 = regVec_1672;
      end
      12'b011010001001 : begin
        _zz__zz_regVec_0 = regVec_1673;
      end
      12'b011010001010 : begin
        _zz__zz_regVec_0 = regVec_1674;
      end
      12'b011010001011 : begin
        _zz__zz_regVec_0 = regVec_1675;
      end
      12'b011010001100 : begin
        _zz__zz_regVec_0 = regVec_1676;
      end
      12'b011010001101 : begin
        _zz__zz_regVec_0 = regVec_1677;
      end
      12'b011010001110 : begin
        _zz__zz_regVec_0 = regVec_1678;
      end
      12'b011010001111 : begin
        _zz__zz_regVec_0 = regVec_1679;
      end
      12'b011010010000 : begin
        _zz__zz_regVec_0 = regVec_1680;
      end
      12'b011010010001 : begin
        _zz__zz_regVec_0 = regVec_1681;
      end
      12'b011010010010 : begin
        _zz__zz_regVec_0 = regVec_1682;
      end
      12'b011010010011 : begin
        _zz__zz_regVec_0 = regVec_1683;
      end
      12'b011010010100 : begin
        _zz__zz_regVec_0 = regVec_1684;
      end
      12'b011010010101 : begin
        _zz__zz_regVec_0 = regVec_1685;
      end
      12'b011010010110 : begin
        _zz__zz_regVec_0 = regVec_1686;
      end
      12'b011010010111 : begin
        _zz__zz_regVec_0 = regVec_1687;
      end
      12'b011010011000 : begin
        _zz__zz_regVec_0 = regVec_1688;
      end
      12'b011010011001 : begin
        _zz__zz_regVec_0 = regVec_1689;
      end
      12'b011010011010 : begin
        _zz__zz_regVec_0 = regVec_1690;
      end
      12'b011010011011 : begin
        _zz__zz_regVec_0 = regVec_1691;
      end
      12'b011010011100 : begin
        _zz__zz_regVec_0 = regVec_1692;
      end
      12'b011010011101 : begin
        _zz__zz_regVec_0 = regVec_1693;
      end
      12'b011010011110 : begin
        _zz__zz_regVec_0 = regVec_1694;
      end
      12'b011010011111 : begin
        _zz__zz_regVec_0 = regVec_1695;
      end
      12'b011010100000 : begin
        _zz__zz_regVec_0 = regVec_1696;
      end
      12'b011010100001 : begin
        _zz__zz_regVec_0 = regVec_1697;
      end
      12'b011010100010 : begin
        _zz__zz_regVec_0 = regVec_1698;
      end
      12'b011010100011 : begin
        _zz__zz_regVec_0 = regVec_1699;
      end
      12'b011010100100 : begin
        _zz__zz_regVec_0 = regVec_1700;
      end
      12'b011010100101 : begin
        _zz__zz_regVec_0 = regVec_1701;
      end
      12'b011010100110 : begin
        _zz__zz_regVec_0 = regVec_1702;
      end
      12'b011010100111 : begin
        _zz__zz_regVec_0 = regVec_1703;
      end
      12'b011010101000 : begin
        _zz__zz_regVec_0 = regVec_1704;
      end
      12'b011010101001 : begin
        _zz__zz_regVec_0 = regVec_1705;
      end
      12'b011010101010 : begin
        _zz__zz_regVec_0 = regVec_1706;
      end
      12'b011010101011 : begin
        _zz__zz_regVec_0 = regVec_1707;
      end
      12'b011010101100 : begin
        _zz__zz_regVec_0 = regVec_1708;
      end
      12'b011010101101 : begin
        _zz__zz_regVec_0 = regVec_1709;
      end
      12'b011010101110 : begin
        _zz__zz_regVec_0 = regVec_1710;
      end
      12'b011010101111 : begin
        _zz__zz_regVec_0 = regVec_1711;
      end
      12'b011010110000 : begin
        _zz__zz_regVec_0 = regVec_1712;
      end
      12'b011010110001 : begin
        _zz__zz_regVec_0 = regVec_1713;
      end
      12'b011010110010 : begin
        _zz__zz_regVec_0 = regVec_1714;
      end
      12'b011010110011 : begin
        _zz__zz_regVec_0 = regVec_1715;
      end
      12'b011010110100 : begin
        _zz__zz_regVec_0 = regVec_1716;
      end
      12'b011010110101 : begin
        _zz__zz_regVec_0 = regVec_1717;
      end
      12'b011010110110 : begin
        _zz__zz_regVec_0 = regVec_1718;
      end
      12'b011010110111 : begin
        _zz__zz_regVec_0 = regVec_1719;
      end
      12'b011010111000 : begin
        _zz__zz_regVec_0 = regVec_1720;
      end
      12'b011010111001 : begin
        _zz__zz_regVec_0 = regVec_1721;
      end
      12'b011010111010 : begin
        _zz__zz_regVec_0 = regVec_1722;
      end
      12'b011010111011 : begin
        _zz__zz_regVec_0 = regVec_1723;
      end
      12'b011010111100 : begin
        _zz__zz_regVec_0 = regVec_1724;
      end
      12'b011010111101 : begin
        _zz__zz_regVec_0 = regVec_1725;
      end
      12'b011010111110 : begin
        _zz__zz_regVec_0 = regVec_1726;
      end
      12'b011010111111 : begin
        _zz__zz_regVec_0 = regVec_1727;
      end
      12'b011011000000 : begin
        _zz__zz_regVec_0 = regVec_1728;
      end
      12'b011011000001 : begin
        _zz__zz_regVec_0 = regVec_1729;
      end
      12'b011011000010 : begin
        _zz__zz_regVec_0 = regVec_1730;
      end
      12'b011011000011 : begin
        _zz__zz_regVec_0 = regVec_1731;
      end
      12'b011011000100 : begin
        _zz__zz_regVec_0 = regVec_1732;
      end
      12'b011011000101 : begin
        _zz__zz_regVec_0 = regVec_1733;
      end
      12'b011011000110 : begin
        _zz__zz_regVec_0 = regVec_1734;
      end
      12'b011011000111 : begin
        _zz__zz_regVec_0 = regVec_1735;
      end
      12'b011011001000 : begin
        _zz__zz_regVec_0 = regVec_1736;
      end
      12'b011011001001 : begin
        _zz__zz_regVec_0 = regVec_1737;
      end
      12'b011011001010 : begin
        _zz__zz_regVec_0 = regVec_1738;
      end
      12'b011011001011 : begin
        _zz__zz_regVec_0 = regVec_1739;
      end
      12'b011011001100 : begin
        _zz__zz_regVec_0 = regVec_1740;
      end
      12'b011011001101 : begin
        _zz__zz_regVec_0 = regVec_1741;
      end
      12'b011011001110 : begin
        _zz__zz_regVec_0 = regVec_1742;
      end
      12'b011011001111 : begin
        _zz__zz_regVec_0 = regVec_1743;
      end
      12'b011011010000 : begin
        _zz__zz_regVec_0 = regVec_1744;
      end
      12'b011011010001 : begin
        _zz__zz_regVec_0 = regVec_1745;
      end
      12'b011011010010 : begin
        _zz__zz_regVec_0 = regVec_1746;
      end
      12'b011011010011 : begin
        _zz__zz_regVec_0 = regVec_1747;
      end
      12'b011011010100 : begin
        _zz__zz_regVec_0 = regVec_1748;
      end
      12'b011011010101 : begin
        _zz__zz_regVec_0 = regVec_1749;
      end
      12'b011011010110 : begin
        _zz__zz_regVec_0 = regVec_1750;
      end
      12'b011011010111 : begin
        _zz__zz_regVec_0 = regVec_1751;
      end
      12'b011011011000 : begin
        _zz__zz_regVec_0 = regVec_1752;
      end
      12'b011011011001 : begin
        _zz__zz_regVec_0 = regVec_1753;
      end
      12'b011011011010 : begin
        _zz__zz_regVec_0 = regVec_1754;
      end
      12'b011011011011 : begin
        _zz__zz_regVec_0 = regVec_1755;
      end
      12'b011011011100 : begin
        _zz__zz_regVec_0 = regVec_1756;
      end
      12'b011011011101 : begin
        _zz__zz_regVec_0 = regVec_1757;
      end
      12'b011011011110 : begin
        _zz__zz_regVec_0 = regVec_1758;
      end
      12'b011011011111 : begin
        _zz__zz_regVec_0 = regVec_1759;
      end
      12'b011011100000 : begin
        _zz__zz_regVec_0 = regVec_1760;
      end
      12'b011011100001 : begin
        _zz__zz_regVec_0 = regVec_1761;
      end
      12'b011011100010 : begin
        _zz__zz_regVec_0 = regVec_1762;
      end
      12'b011011100011 : begin
        _zz__zz_regVec_0 = regVec_1763;
      end
      12'b011011100100 : begin
        _zz__zz_regVec_0 = regVec_1764;
      end
      12'b011011100101 : begin
        _zz__zz_regVec_0 = regVec_1765;
      end
      12'b011011100110 : begin
        _zz__zz_regVec_0 = regVec_1766;
      end
      12'b011011100111 : begin
        _zz__zz_regVec_0 = regVec_1767;
      end
      12'b011011101000 : begin
        _zz__zz_regVec_0 = regVec_1768;
      end
      12'b011011101001 : begin
        _zz__zz_regVec_0 = regVec_1769;
      end
      12'b011011101010 : begin
        _zz__zz_regVec_0 = regVec_1770;
      end
      12'b011011101011 : begin
        _zz__zz_regVec_0 = regVec_1771;
      end
      12'b011011101100 : begin
        _zz__zz_regVec_0 = regVec_1772;
      end
      12'b011011101101 : begin
        _zz__zz_regVec_0 = regVec_1773;
      end
      12'b011011101110 : begin
        _zz__zz_regVec_0 = regVec_1774;
      end
      12'b011011101111 : begin
        _zz__zz_regVec_0 = regVec_1775;
      end
      12'b011011110000 : begin
        _zz__zz_regVec_0 = regVec_1776;
      end
      12'b011011110001 : begin
        _zz__zz_regVec_0 = regVec_1777;
      end
      12'b011011110010 : begin
        _zz__zz_regVec_0 = regVec_1778;
      end
      12'b011011110011 : begin
        _zz__zz_regVec_0 = regVec_1779;
      end
      12'b011011110100 : begin
        _zz__zz_regVec_0 = regVec_1780;
      end
      12'b011011110101 : begin
        _zz__zz_regVec_0 = regVec_1781;
      end
      12'b011011110110 : begin
        _zz__zz_regVec_0 = regVec_1782;
      end
      12'b011011110111 : begin
        _zz__zz_regVec_0 = regVec_1783;
      end
      12'b011011111000 : begin
        _zz__zz_regVec_0 = regVec_1784;
      end
      12'b011011111001 : begin
        _zz__zz_regVec_0 = regVec_1785;
      end
      12'b011011111010 : begin
        _zz__zz_regVec_0 = regVec_1786;
      end
      12'b011011111011 : begin
        _zz__zz_regVec_0 = regVec_1787;
      end
      12'b011011111100 : begin
        _zz__zz_regVec_0 = regVec_1788;
      end
      12'b011011111101 : begin
        _zz__zz_regVec_0 = regVec_1789;
      end
      12'b011011111110 : begin
        _zz__zz_regVec_0 = regVec_1790;
      end
      12'b011011111111 : begin
        _zz__zz_regVec_0 = regVec_1791;
      end
      12'b011100000000 : begin
        _zz__zz_regVec_0 = regVec_1792;
      end
      12'b011100000001 : begin
        _zz__zz_regVec_0 = regVec_1793;
      end
      12'b011100000010 : begin
        _zz__zz_regVec_0 = regVec_1794;
      end
      12'b011100000011 : begin
        _zz__zz_regVec_0 = regVec_1795;
      end
      12'b011100000100 : begin
        _zz__zz_regVec_0 = regVec_1796;
      end
      12'b011100000101 : begin
        _zz__zz_regVec_0 = regVec_1797;
      end
      12'b011100000110 : begin
        _zz__zz_regVec_0 = regVec_1798;
      end
      12'b011100000111 : begin
        _zz__zz_regVec_0 = regVec_1799;
      end
      12'b011100001000 : begin
        _zz__zz_regVec_0 = regVec_1800;
      end
      12'b011100001001 : begin
        _zz__zz_regVec_0 = regVec_1801;
      end
      12'b011100001010 : begin
        _zz__zz_regVec_0 = regVec_1802;
      end
      12'b011100001011 : begin
        _zz__zz_regVec_0 = regVec_1803;
      end
      12'b011100001100 : begin
        _zz__zz_regVec_0 = regVec_1804;
      end
      12'b011100001101 : begin
        _zz__zz_regVec_0 = regVec_1805;
      end
      12'b011100001110 : begin
        _zz__zz_regVec_0 = regVec_1806;
      end
      12'b011100001111 : begin
        _zz__zz_regVec_0 = regVec_1807;
      end
      12'b011100010000 : begin
        _zz__zz_regVec_0 = regVec_1808;
      end
      12'b011100010001 : begin
        _zz__zz_regVec_0 = regVec_1809;
      end
      12'b011100010010 : begin
        _zz__zz_regVec_0 = regVec_1810;
      end
      12'b011100010011 : begin
        _zz__zz_regVec_0 = regVec_1811;
      end
      12'b011100010100 : begin
        _zz__zz_regVec_0 = regVec_1812;
      end
      12'b011100010101 : begin
        _zz__zz_regVec_0 = regVec_1813;
      end
      12'b011100010110 : begin
        _zz__zz_regVec_0 = regVec_1814;
      end
      12'b011100010111 : begin
        _zz__zz_regVec_0 = regVec_1815;
      end
      12'b011100011000 : begin
        _zz__zz_regVec_0 = regVec_1816;
      end
      12'b011100011001 : begin
        _zz__zz_regVec_0 = regVec_1817;
      end
      12'b011100011010 : begin
        _zz__zz_regVec_0 = regVec_1818;
      end
      12'b011100011011 : begin
        _zz__zz_regVec_0 = regVec_1819;
      end
      12'b011100011100 : begin
        _zz__zz_regVec_0 = regVec_1820;
      end
      12'b011100011101 : begin
        _zz__zz_regVec_0 = regVec_1821;
      end
      12'b011100011110 : begin
        _zz__zz_regVec_0 = regVec_1822;
      end
      12'b011100011111 : begin
        _zz__zz_regVec_0 = regVec_1823;
      end
      12'b011100100000 : begin
        _zz__zz_regVec_0 = regVec_1824;
      end
      12'b011100100001 : begin
        _zz__zz_regVec_0 = regVec_1825;
      end
      12'b011100100010 : begin
        _zz__zz_regVec_0 = regVec_1826;
      end
      12'b011100100011 : begin
        _zz__zz_regVec_0 = regVec_1827;
      end
      12'b011100100100 : begin
        _zz__zz_regVec_0 = regVec_1828;
      end
      12'b011100100101 : begin
        _zz__zz_regVec_0 = regVec_1829;
      end
      12'b011100100110 : begin
        _zz__zz_regVec_0 = regVec_1830;
      end
      12'b011100100111 : begin
        _zz__zz_regVec_0 = regVec_1831;
      end
      12'b011100101000 : begin
        _zz__zz_regVec_0 = regVec_1832;
      end
      12'b011100101001 : begin
        _zz__zz_regVec_0 = regVec_1833;
      end
      12'b011100101010 : begin
        _zz__zz_regVec_0 = regVec_1834;
      end
      12'b011100101011 : begin
        _zz__zz_regVec_0 = regVec_1835;
      end
      12'b011100101100 : begin
        _zz__zz_regVec_0 = regVec_1836;
      end
      12'b011100101101 : begin
        _zz__zz_regVec_0 = regVec_1837;
      end
      12'b011100101110 : begin
        _zz__zz_regVec_0 = regVec_1838;
      end
      12'b011100101111 : begin
        _zz__zz_regVec_0 = regVec_1839;
      end
      12'b011100110000 : begin
        _zz__zz_regVec_0 = regVec_1840;
      end
      12'b011100110001 : begin
        _zz__zz_regVec_0 = regVec_1841;
      end
      12'b011100110010 : begin
        _zz__zz_regVec_0 = regVec_1842;
      end
      12'b011100110011 : begin
        _zz__zz_regVec_0 = regVec_1843;
      end
      12'b011100110100 : begin
        _zz__zz_regVec_0 = regVec_1844;
      end
      12'b011100110101 : begin
        _zz__zz_regVec_0 = regVec_1845;
      end
      12'b011100110110 : begin
        _zz__zz_regVec_0 = regVec_1846;
      end
      12'b011100110111 : begin
        _zz__zz_regVec_0 = regVec_1847;
      end
      12'b011100111000 : begin
        _zz__zz_regVec_0 = regVec_1848;
      end
      12'b011100111001 : begin
        _zz__zz_regVec_0 = regVec_1849;
      end
      12'b011100111010 : begin
        _zz__zz_regVec_0 = regVec_1850;
      end
      12'b011100111011 : begin
        _zz__zz_regVec_0 = regVec_1851;
      end
      12'b011100111100 : begin
        _zz__zz_regVec_0 = regVec_1852;
      end
      12'b011100111101 : begin
        _zz__zz_regVec_0 = regVec_1853;
      end
      12'b011100111110 : begin
        _zz__zz_regVec_0 = regVec_1854;
      end
      12'b011100111111 : begin
        _zz__zz_regVec_0 = regVec_1855;
      end
      12'b011101000000 : begin
        _zz__zz_regVec_0 = regVec_1856;
      end
      12'b011101000001 : begin
        _zz__zz_regVec_0 = regVec_1857;
      end
      12'b011101000010 : begin
        _zz__zz_regVec_0 = regVec_1858;
      end
      12'b011101000011 : begin
        _zz__zz_regVec_0 = regVec_1859;
      end
      12'b011101000100 : begin
        _zz__zz_regVec_0 = regVec_1860;
      end
      12'b011101000101 : begin
        _zz__zz_regVec_0 = regVec_1861;
      end
      12'b011101000110 : begin
        _zz__zz_regVec_0 = regVec_1862;
      end
      12'b011101000111 : begin
        _zz__zz_regVec_0 = regVec_1863;
      end
      12'b011101001000 : begin
        _zz__zz_regVec_0 = regVec_1864;
      end
      12'b011101001001 : begin
        _zz__zz_regVec_0 = regVec_1865;
      end
      12'b011101001010 : begin
        _zz__zz_regVec_0 = regVec_1866;
      end
      12'b011101001011 : begin
        _zz__zz_regVec_0 = regVec_1867;
      end
      12'b011101001100 : begin
        _zz__zz_regVec_0 = regVec_1868;
      end
      12'b011101001101 : begin
        _zz__zz_regVec_0 = regVec_1869;
      end
      12'b011101001110 : begin
        _zz__zz_regVec_0 = regVec_1870;
      end
      12'b011101001111 : begin
        _zz__zz_regVec_0 = regVec_1871;
      end
      12'b011101010000 : begin
        _zz__zz_regVec_0 = regVec_1872;
      end
      12'b011101010001 : begin
        _zz__zz_regVec_0 = regVec_1873;
      end
      12'b011101010010 : begin
        _zz__zz_regVec_0 = regVec_1874;
      end
      12'b011101010011 : begin
        _zz__zz_regVec_0 = regVec_1875;
      end
      12'b011101010100 : begin
        _zz__zz_regVec_0 = regVec_1876;
      end
      12'b011101010101 : begin
        _zz__zz_regVec_0 = regVec_1877;
      end
      12'b011101010110 : begin
        _zz__zz_regVec_0 = regVec_1878;
      end
      12'b011101010111 : begin
        _zz__zz_regVec_0 = regVec_1879;
      end
      12'b011101011000 : begin
        _zz__zz_regVec_0 = regVec_1880;
      end
      12'b011101011001 : begin
        _zz__zz_regVec_0 = regVec_1881;
      end
      12'b011101011010 : begin
        _zz__zz_regVec_0 = regVec_1882;
      end
      12'b011101011011 : begin
        _zz__zz_regVec_0 = regVec_1883;
      end
      12'b011101011100 : begin
        _zz__zz_regVec_0 = regVec_1884;
      end
      12'b011101011101 : begin
        _zz__zz_regVec_0 = regVec_1885;
      end
      12'b011101011110 : begin
        _zz__zz_regVec_0 = regVec_1886;
      end
      12'b011101011111 : begin
        _zz__zz_regVec_0 = regVec_1887;
      end
      12'b011101100000 : begin
        _zz__zz_regVec_0 = regVec_1888;
      end
      12'b011101100001 : begin
        _zz__zz_regVec_0 = regVec_1889;
      end
      12'b011101100010 : begin
        _zz__zz_regVec_0 = regVec_1890;
      end
      12'b011101100011 : begin
        _zz__zz_regVec_0 = regVec_1891;
      end
      12'b011101100100 : begin
        _zz__zz_regVec_0 = regVec_1892;
      end
      12'b011101100101 : begin
        _zz__zz_regVec_0 = regVec_1893;
      end
      12'b011101100110 : begin
        _zz__zz_regVec_0 = regVec_1894;
      end
      12'b011101100111 : begin
        _zz__zz_regVec_0 = regVec_1895;
      end
      12'b011101101000 : begin
        _zz__zz_regVec_0 = regVec_1896;
      end
      12'b011101101001 : begin
        _zz__zz_regVec_0 = regVec_1897;
      end
      12'b011101101010 : begin
        _zz__zz_regVec_0 = regVec_1898;
      end
      12'b011101101011 : begin
        _zz__zz_regVec_0 = regVec_1899;
      end
      12'b011101101100 : begin
        _zz__zz_regVec_0 = regVec_1900;
      end
      12'b011101101101 : begin
        _zz__zz_regVec_0 = regVec_1901;
      end
      12'b011101101110 : begin
        _zz__zz_regVec_0 = regVec_1902;
      end
      12'b011101101111 : begin
        _zz__zz_regVec_0 = regVec_1903;
      end
      12'b011101110000 : begin
        _zz__zz_regVec_0 = regVec_1904;
      end
      12'b011101110001 : begin
        _zz__zz_regVec_0 = regVec_1905;
      end
      12'b011101110010 : begin
        _zz__zz_regVec_0 = regVec_1906;
      end
      12'b011101110011 : begin
        _zz__zz_regVec_0 = regVec_1907;
      end
      12'b011101110100 : begin
        _zz__zz_regVec_0 = regVec_1908;
      end
      12'b011101110101 : begin
        _zz__zz_regVec_0 = regVec_1909;
      end
      12'b011101110110 : begin
        _zz__zz_regVec_0 = regVec_1910;
      end
      12'b011101110111 : begin
        _zz__zz_regVec_0 = regVec_1911;
      end
      12'b011101111000 : begin
        _zz__zz_regVec_0 = regVec_1912;
      end
      12'b011101111001 : begin
        _zz__zz_regVec_0 = regVec_1913;
      end
      12'b011101111010 : begin
        _zz__zz_regVec_0 = regVec_1914;
      end
      12'b011101111011 : begin
        _zz__zz_regVec_0 = regVec_1915;
      end
      12'b011101111100 : begin
        _zz__zz_regVec_0 = regVec_1916;
      end
      12'b011101111101 : begin
        _zz__zz_regVec_0 = regVec_1917;
      end
      12'b011101111110 : begin
        _zz__zz_regVec_0 = regVec_1918;
      end
      12'b011101111111 : begin
        _zz__zz_regVec_0 = regVec_1919;
      end
      12'b011110000000 : begin
        _zz__zz_regVec_0 = regVec_1920;
      end
      12'b011110000001 : begin
        _zz__zz_regVec_0 = regVec_1921;
      end
      12'b011110000010 : begin
        _zz__zz_regVec_0 = regVec_1922;
      end
      12'b011110000011 : begin
        _zz__zz_regVec_0 = regVec_1923;
      end
      12'b011110000100 : begin
        _zz__zz_regVec_0 = regVec_1924;
      end
      12'b011110000101 : begin
        _zz__zz_regVec_0 = regVec_1925;
      end
      12'b011110000110 : begin
        _zz__zz_regVec_0 = regVec_1926;
      end
      12'b011110000111 : begin
        _zz__zz_regVec_0 = regVec_1927;
      end
      12'b011110001000 : begin
        _zz__zz_regVec_0 = regVec_1928;
      end
      12'b011110001001 : begin
        _zz__zz_regVec_0 = regVec_1929;
      end
      12'b011110001010 : begin
        _zz__zz_regVec_0 = regVec_1930;
      end
      12'b011110001011 : begin
        _zz__zz_regVec_0 = regVec_1931;
      end
      12'b011110001100 : begin
        _zz__zz_regVec_0 = regVec_1932;
      end
      12'b011110001101 : begin
        _zz__zz_regVec_0 = regVec_1933;
      end
      12'b011110001110 : begin
        _zz__zz_regVec_0 = regVec_1934;
      end
      12'b011110001111 : begin
        _zz__zz_regVec_0 = regVec_1935;
      end
      12'b011110010000 : begin
        _zz__zz_regVec_0 = regVec_1936;
      end
      12'b011110010001 : begin
        _zz__zz_regVec_0 = regVec_1937;
      end
      12'b011110010010 : begin
        _zz__zz_regVec_0 = regVec_1938;
      end
      12'b011110010011 : begin
        _zz__zz_regVec_0 = regVec_1939;
      end
      12'b011110010100 : begin
        _zz__zz_regVec_0 = regVec_1940;
      end
      12'b011110010101 : begin
        _zz__zz_regVec_0 = regVec_1941;
      end
      12'b011110010110 : begin
        _zz__zz_regVec_0 = regVec_1942;
      end
      12'b011110010111 : begin
        _zz__zz_regVec_0 = regVec_1943;
      end
      12'b011110011000 : begin
        _zz__zz_regVec_0 = regVec_1944;
      end
      12'b011110011001 : begin
        _zz__zz_regVec_0 = regVec_1945;
      end
      12'b011110011010 : begin
        _zz__zz_regVec_0 = regVec_1946;
      end
      12'b011110011011 : begin
        _zz__zz_regVec_0 = regVec_1947;
      end
      12'b011110011100 : begin
        _zz__zz_regVec_0 = regVec_1948;
      end
      12'b011110011101 : begin
        _zz__zz_regVec_0 = regVec_1949;
      end
      12'b011110011110 : begin
        _zz__zz_regVec_0 = regVec_1950;
      end
      12'b011110011111 : begin
        _zz__zz_regVec_0 = regVec_1951;
      end
      12'b011110100000 : begin
        _zz__zz_regVec_0 = regVec_1952;
      end
      12'b011110100001 : begin
        _zz__zz_regVec_0 = regVec_1953;
      end
      12'b011110100010 : begin
        _zz__zz_regVec_0 = regVec_1954;
      end
      12'b011110100011 : begin
        _zz__zz_regVec_0 = regVec_1955;
      end
      12'b011110100100 : begin
        _zz__zz_regVec_0 = regVec_1956;
      end
      12'b011110100101 : begin
        _zz__zz_regVec_0 = regVec_1957;
      end
      12'b011110100110 : begin
        _zz__zz_regVec_0 = regVec_1958;
      end
      12'b011110100111 : begin
        _zz__zz_regVec_0 = regVec_1959;
      end
      12'b011110101000 : begin
        _zz__zz_regVec_0 = regVec_1960;
      end
      12'b011110101001 : begin
        _zz__zz_regVec_0 = regVec_1961;
      end
      12'b011110101010 : begin
        _zz__zz_regVec_0 = regVec_1962;
      end
      12'b011110101011 : begin
        _zz__zz_regVec_0 = regVec_1963;
      end
      12'b011110101100 : begin
        _zz__zz_regVec_0 = regVec_1964;
      end
      12'b011110101101 : begin
        _zz__zz_regVec_0 = regVec_1965;
      end
      12'b011110101110 : begin
        _zz__zz_regVec_0 = regVec_1966;
      end
      12'b011110101111 : begin
        _zz__zz_regVec_0 = regVec_1967;
      end
      12'b011110110000 : begin
        _zz__zz_regVec_0 = regVec_1968;
      end
      12'b011110110001 : begin
        _zz__zz_regVec_0 = regVec_1969;
      end
      12'b011110110010 : begin
        _zz__zz_regVec_0 = regVec_1970;
      end
      12'b011110110011 : begin
        _zz__zz_regVec_0 = regVec_1971;
      end
      12'b011110110100 : begin
        _zz__zz_regVec_0 = regVec_1972;
      end
      12'b011110110101 : begin
        _zz__zz_regVec_0 = regVec_1973;
      end
      12'b011110110110 : begin
        _zz__zz_regVec_0 = regVec_1974;
      end
      12'b011110110111 : begin
        _zz__zz_regVec_0 = regVec_1975;
      end
      12'b011110111000 : begin
        _zz__zz_regVec_0 = regVec_1976;
      end
      12'b011110111001 : begin
        _zz__zz_regVec_0 = regVec_1977;
      end
      12'b011110111010 : begin
        _zz__zz_regVec_0 = regVec_1978;
      end
      12'b011110111011 : begin
        _zz__zz_regVec_0 = regVec_1979;
      end
      12'b011110111100 : begin
        _zz__zz_regVec_0 = regVec_1980;
      end
      12'b011110111101 : begin
        _zz__zz_regVec_0 = regVec_1981;
      end
      12'b011110111110 : begin
        _zz__zz_regVec_0 = regVec_1982;
      end
      12'b011110111111 : begin
        _zz__zz_regVec_0 = regVec_1983;
      end
      12'b011111000000 : begin
        _zz__zz_regVec_0 = regVec_1984;
      end
      12'b011111000001 : begin
        _zz__zz_regVec_0 = regVec_1985;
      end
      12'b011111000010 : begin
        _zz__zz_regVec_0 = regVec_1986;
      end
      12'b011111000011 : begin
        _zz__zz_regVec_0 = regVec_1987;
      end
      12'b011111000100 : begin
        _zz__zz_regVec_0 = regVec_1988;
      end
      12'b011111000101 : begin
        _zz__zz_regVec_0 = regVec_1989;
      end
      12'b011111000110 : begin
        _zz__zz_regVec_0 = regVec_1990;
      end
      12'b011111000111 : begin
        _zz__zz_regVec_0 = regVec_1991;
      end
      12'b011111001000 : begin
        _zz__zz_regVec_0 = regVec_1992;
      end
      12'b011111001001 : begin
        _zz__zz_regVec_0 = regVec_1993;
      end
      12'b011111001010 : begin
        _zz__zz_regVec_0 = regVec_1994;
      end
      12'b011111001011 : begin
        _zz__zz_regVec_0 = regVec_1995;
      end
      12'b011111001100 : begin
        _zz__zz_regVec_0 = regVec_1996;
      end
      12'b011111001101 : begin
        _zz__zz_regVec_0 = regVec_1997;
      end
      12'b011111001110 : begin
        _zz__zz_regVec_0 = regVec_1998;
      end
      12'b011111001111 : begin
        _zz__zz_regVec_0 = regVec_1999;
      end
      12'b011111010000 : begin
        _zz__zz_regVec_0 = regVec_2000;
      end
      12'b011111010001 : begin
        _zz__zz_regVec_0 = regVec_2001;
      end
      12'b011111010010 : begin
        _zz__zz_regVec_0 = regVec_2002;
      end
      12'b011111010011 : begin
        _zz__zz_regVec_0 = regVec_2003;
      end
      12'b011111010100 : begin
        _zz__zz_regVec_0 = regVec_2004;
      end
      12'b011111010101 : begin
        _zz__zz_regVec_0 = regVec_2005;
      end
      12'b011111010110 : begin
        _zz__zz_regVec_0 = regVec_2006;
      end
      12'b011111010111 : begin
        _zz__zz_regVec_0 = regVec_2007;
      end
      12'b011111011000 : begin
        _zz__zz_regVec_0 = regVec_2008;
      end
      12'b011111011001 : begin
        _zz__zz_regVec_0 = regVec_2009;
      end
      12'b011111011010 : begin
        _zz__zz_regVec_0 = regVec_2010;
      end
      12'b011111011011 : begin
        _zz__zz_regVec_0 = regVec_2011;
      end
      12'b011111011100 : begin
        _zz__zz_regVec_0 = regVec_2012;
      end
      12'b011111011101 : begin
        _zz__zz_regVec_0 = regVec_2013;
      end
      12'b011111011110 : begin
        _zz__zz_regVec_0 = regVec_2014;
      end
      12'b011111011111 : begin
        _zz__zz_regVec_0 = regVec_2015;
      end
      12'b011111100000 : begin
        _zz__zz_regVec_0 = regVec_2016;
      end
      12'b011111100001 : begin
        _zz__zz_regVec_0 = regVec_2017;
      end
      12'b011111100010 : begin
        _zz__zz_regVec_0 = regVec_2018;
      end
      12'b011111100011 : begin
        _zz__zz_regVec_0 = regVec_2019;
      end
      12'b011111100100 : begin
        _zz__zz_regVec_0 = regVec_2020;
      end
      12'b011111100101 : begin
        _zz__zz_regVec_0 = regVec_2021;
      end
      12'b011111100110 : begin
        _zz__zz_regVec_0 = regVec_2022;
      end
      12'b011111100111 : begin
        _zz__zz_regVec_0 = regVec_2023;
      end
      12'b011111101000 : begin
        _zz__zz_regVec_0 = regVec_2024;
      end
      12'b011111101001 : begin
        _zz__zz_regVec_0 = regVec_2025;
      end
      12'b011111101010 : begin
        _zz__zz_regVec_0 = regVec_2026;
      end
      12'b011111101011 : begin
        _zz__zz_regVec_0 = regVec_2027;
      end
      12'b011111101100 : begin
        _zz__zz_regVec_0 = regVec_2028;
      end
      12'b011111101101 : begin
        _zz__zz_regVec_0 = regVec_2029;
      end
      12'b011111101110 : begin
        _zz__zz_regVec_0 = regVec_2030;
      end
      12'b011111101111 : begin
        _zz__zz_regVec_0 = regVec_2031;
      end
      12'b011111110000 : begin
        _zz__zz_regVec_0 = regVec_2032;
      end
      12'b011111110001 : begin
        _zz__zz_regVec_0 = regVec_2033;
      end
      12'b011111110010 : begin
        _zz__zz_regVec_0 = regVec_2034;
      end
      12'b011111110011 : begin
        _zz__zz_regVec_0 = regVec_2035;
      end
      12'b011111110100 : begin
        _zz__zz_regVec_0 = regVec_2036;
      end
      12'b011111110101 : begin
        _zz__zz_regVec_0 = regVec_2037;
      end
      12'b011111110110 : begin
        _zz__zz_regVec_0 = regVec_2038;
      end
      12'b011111110111 : begin
        _zz__zz_regVec_0 = regVec_2039;
      end
      12'b011111111000 : begin
        _zz__zz_regVec_0 = regVec_2040;
      end
      12'b011111111001 : begin
        _zz__zz_regVec_0 = regVec_2041;
      end
      12'b011111111010 : begin
        _zz__zz_regVec_0 = regVec_2042;
      end
      12'b011111111011 : begin
        _zz__zz_regVec_0 = regVec_2043;
      end
      12'b011111111100 : begin
        _zz__zz_regVec_0 = regVec_2044;
      end
      12'b011111111101 : begin
        _zz__zz_regVec_0 = regVec_2045;
      end
      12'b011111111110 : begin
        _zz__zz_regVec_0 = regVec_2046;
      end
      12'b011111111111 : begin
        _zz__zz_regVec_0 = regVec_2047;
      end
      12'b100000000000 : begin
        _zz__zz_regVec_0 = regVec_2048;
      end
      12'b100000000001 : begin
        _zz__zz_regVec_0 = regVec_2049;
      end
      12'b100000000010 : begin
        _zz__zz_regVec_0 = regVec_2050;
      end
      12'b100000000011 : begin
        _zz__zz_regVec_0 = regVec_2051;
      end
      12'b100000000100 : begin
        _zz__zz_regVec_0 = regVec_2052;
      end
      12'b100000000101 : begin
        _zz__zz_regVec_0 = regVec_2053;
      end
      12'b100000000110 : begin
        _zz__zz_regVec_0 = regVec_2054;
      end
      12'b100000000111 : begin
        _zz__zz_regVec_0 = regVec_2055;
      end
      12'b100000001000 : begin
        _zz__zz_regVec_0 = regVec_2056;
      end
      12'b100000001001 : begin
        _zz__zz_regVec_0 = regVec_2057;
      end
      12'b100000001010 : begin
        _zz__zz_regVec_0 = regVec_2058;
      end
      12'b100000001011 : begin
        _zz__zz_regVec_0 = regVec_2059;
      end
      12'b100000001100 : begin
        _zz__zz_regVec_0 = regVec_2060;
      end
      12'b100000001101 : begin
        _zz__zz_regVec_0 = regVec_2061;
      end
      12'b100000001110 : begin
        _zz__zz_regVec_0 = regVec_2062;
      end
      12'b100000001111 : begin
        _zz__zz_regVec_0 = regVec_2063;
      end
      12'b100000010000 : begin
        _zz__zz_regVec_0 = regVec_2064;
      end
      12'b100000010001 : begin
        _zz__zz_regVec_0 = regVec_2065;
      end
      12'b100000010010 : begin
        _zz__zz_regVec_0 = regVec_2066;
      end
      12'b100000010011 : begin
        _zz__zz_regVec_0 = regVec_2067;
      end
      12'b100000010100 : begin
        _zz__zz_regVec_0 = regVec_2068;
      end
      12'b100000010101 : begin
        _zz__zz_regVec_0 = regVec_2069;
      end
      12'b100000010110 : begin
        _zz__zz_regVec_0 = regVec_2070;
      end
      12'b100000010111 : begin
        _zz__zz_regVec_0 = regVec_2071;
      end
      12'b100000011000 : begin
        _zz__zz_regVec_0 = regVec_2072;
      end
      12'b100000011001 : begin
        _zz__zz_regVec_0 = regVec_2073;
      end
      12'b100000011010 : begin
        _zz__zz_regVec_0 = regVec_2074;
      end
      12'b100000011011 : begin
        _zz__zz_regVec_0 = regVec_2075;
      end
      12'b100000011100 : begin
        _zz__zz_regVec_0 = regVec_2076;
      end
      12'b100000011101 : begin
        _zz__zz_regVec_0 = regVec_2077;
      end
      12'b100000011110 : begin
        _zz__zz_regVec_0 = regVec_2078;
      end
      12'b100000011111 : begin
        _zz__zz_regVec_0 = regVec_2079;
      end
      12'b100000100000 : begin
        _zz__zz_regVec_0 = regVec_2080;
      end
      12'b100000100001 : begin
        _zz__zz_regVec_0 = regVec_2081;
      end
      12'b100000100010 : begin
        _zz__zz_regVec_0 = regVec_2082;
      end
      12'b100000100011 : begin
        _zz__zz_regVec_0 = regVec_2083;
      end
      12'b100000100100 : begin
        _zz__zz_regVec_0 = regVec_2084;
      end
      12'b100000100101 : begin
        _zz__zz_regVec_0 = regVec_2085;
      end
      12'b100000100110 : begin
        _zz__zz_regVec_0 = regVec_2086;
      end
      12'b100000100111 : begin
        _zz__zz_regVec_0 = regVec_2087;
      end
      12'b100000101000 : begin
        _zz__zz_regVec_0 = regVec_2088;
      end
      12'b100000101001 : begin
        _zz__zz_regVec_0 = regVec_2089;
      end
      12'b100000101010 : begin
        _zz__zz_regVec_0 = regVec_2090;
      end
      12'b100000101011 : begin
        _zz__zz_regVec_0 = regVec_2091;
      end
      12'b100000101100 : begin
        _zz__zz_regVec_0 = regVec_2092;
      end
      12'b100000101101 : begin
        _zz__zz_regVec_0 = regVec_2093;
      end
      12'b100000101110 : begin
        _zz__zz_regVec_0 = regVec_2094;
      end
      12'b100000101111 : begin
        _zz__zz_regVec_0 = regVec_2095;
      end
      12'b100000110000 : begin
        _zz__zz_regVec_0 = regVec_2096;
      end
      12'b100000110001 : begin
        _zz__zz_regVec_0 = regVec_2097;
      end
      12'b100000110010 : begin
        _zz__zz_regVec_0 = regVec_2098;
      end
      12'b100000110011 : begin
        _zz__zz_regVec_0 = regVec_2099;
      end
      12'b100000110100 : begin
        _zz__zz_regVec_0 = regVec_2100;
      end
      12'b100000110101 : begin
        _zz__zz_regVec_0 = regVec_2101;
      end
      12'b100000110110 : begin
        _zz__zz_regVec_0 = regVec_2102;
      end
      12'b100000110111 : begin
        _zz__zz_regVec_0 = regVec_2103;
      end
      12'b100000111000 : begin
        _zz__zz_regVec_0 = regVec_2104;
      end
      12'b100000111001 : begin
        _zz__zz_regVec_0 = regVec_2105;
      end
      12'b100000111010 : begin
        _zz__zz_regVec_0 = regVec_2106;
      end
      12'b100000111011 : begin
        _zz__zz_regVec_0 = regVec_2107;
      end
      12'b100000111100 : begin
        _zz__zz_regVec_0 = regVec_2108;
      end
      12'b100000111101 : begin
        _zz__zz_regVec_0 = regVec_2109;
      end
      12'b100000111110 : begin
        _zz__zz_regVec_0 = regVec_2110;
      end
      12'b100000111111 : begin
        _zz__zz_regVec_0 = regVec_2111;
      end
      12'b100001000000 : begin
        _zz__zz_regVec_0 = regVec_2112;
      end
      12'b100001000001 : begin
        _zz__zz_regVec_0 = regVec_2113;
      end
      12'b100001000010 : begin
        _zz__zz_regVec_0 = regVec_2114;
      end
      12'b100001000011 : begin
        _zz__zz_regVec_0 = regVec_2115;
      end
      12'b100001000100 : begin
        _zz__zz_regVec_0 = regVec_2116;
      end
      12'b100001000101 : begin
        _zz__zz_regVec_0 = regVec_2117;
      end
      12'b100001000110 : begin
        _zz__zz_regVec_0 = regVec_2118;
      end
      12'b100001000111 : begin
        _zz__zz_regVec_0 = regVec_2119;
      end
      12'b100001001000 : begin
        _zz__zz_regVec_0 = regVec_2120;
      end
      12'b100001001001 : begin
        _zz__zz_regVec_0 = regVec_2121;
      end
      12'b100001001010 : begin
        _zz__zz_regVec_0 = regVec_2122;
      end
      12'b100001001011 : begin
        _zz__zz_regVec_0 = regVec_2123;
      end
      12'b100001001100 : begin
        _zz__zz_regVec_0 = regVec_2124;
      end
      12'b100001001101 : begin
        _zz__zz_regVec_0 = regVec_2125;
      end
      12'b100001001110 : begin
        _zz__zz_regVec_0 = regVec_2126;
      end
      12'b100001001111 : begin
        _zz__zz_regVec_0 = regVec_2127;
      end
      12'b100001010000 : begin
        _zz__zz_regVec_0 = regVec_2128;
      end
      12'b100001010001 : begin
        _zz__zz_regVec_0 = regVec_2129;
      end
      12'b100001010010 : begin
        _zz__zz_regVec_0 = regVec_2130;
      end
      12'b100001010011 : begin
        _zz__zz_regVec_0 = regVec_2131;
      end
      12'b100001010100 : begin
        _zz__zz_regVec_0 = regVec_2132;
      end
      12'b100001010101 : begin
        _zz__zz_regVec_0 = regVec_2133;
      end
      12'b100001010110 : begin
        _zz__zz_regVec_0 = regVec_2134;
      end
      12'b100001010111 : begin
        _zz__zz_regVec_0 = regVec_2135;
      end
      12'b100001011000 : begin
        _zz__zz_regVec_0 = regVec_2136;
      end
      12'b100001011001 : begin
        _zz__zz_regVec_0 = regVec_2137;
      end
      12'b100001011010 : begin
        _zz__zz_regVec_0 = regVec_2138;
      end
      12'b100001011011 : begin
        _zz__zz_regVec_0 = regVec_2139;
      end
      12'b100001011100 : begin
        _zz__zz_regVec_0 = regVec_2140;
      end
      12'b100001011101 : begin
        _zz__zz_regVec_0 = regVec_2141;
      end
      12'b100001011110 : begin
        _zz__zz_regVec_0 = regVec_2142;
      end
      12'b100001011111 : begin
        _zz__zz_regVec_0 = regVec_2143;
      end
      12'b100001100000 : begin
        _zz__zz_regVec_0 = regVec_2144;
      end
      12'b100001100001 : begin
        _zz__zz_regVec_0 = regVec_2145;
      end
      12'b100001100010 : begin
        _zz__zz_regVec_0 = regVec_2146;
      end
      12'b100001100011 : begin
        _zz__zz_regVec_0 = regVec_2147;
      end
      12'b100001100100 : begin
        _zz__zz_regVec_0 = regVec_2148;
      end
      12'b100001100101 : begin
        _zz__zz_regVec_0 = regVec_2149;
      end
      12'b100001100110 : begin
        _zz__zz_regVec_0 = regVec_2150;
      end
      12'b100001100111 : begin
        _zz__zz_regVec_0 = regVec_2151;
      end
      12'b100001101000 : begin
        _zz__zz_regVec_0 = regVec_2152;
      end
      12'b100001101001 : begin
        _zz__zz_regVec_0 = regVec_2153;
      end
      12'b100001101010 : begin
        _zz__zz_regVec_0 = regVec_2154;
      end
      12'b100001101011 : begin
        _zz__zz_regVec_0 = regVec_2155;
      end
      12'b100001101100 : begin
        _zz__zz_regVec_0 = regVec_2156;
      end
      12'b100001101101 : begin
        _zz__zz_regVec_0 = regVec_2157;
      end
      12'b100001101110 : begin
        _zz__zz_regVec_0 = regVec_2158;
      end
      12'b100001101111 : begin
        _zz__zz_regVec_0 = regVec_2159;
      end
      12'b100001110000 : begin
        _zz__zz_regVec_0 = regVec_2160;
      end
      12'b100001110001 : begin
        _zz__zz_regVec_0 = regVec_2161;
      end
      12'b100001110010 : begin
        _zz__zz_regVec_0 = regVec_2162;
      end
      12'b100001110011 : begin
        _zz__zz_regVec_0 = regVec_2163;
      end
      12'b100001110100 : begin
        _zz__zz_regVec_0 = regVec_2164;
      end
      12'b100001110101 : begin
        _zz__zz_regVec_0 = regVec_2165;
      end
      12'b100001110110 : begin
        _zz__zz_regVec_0 = regVec_2166;
      end
      12'b100001110111 : begin
        _zz__zz_regVec_0 = regVec_2167;
      end
      12'b100001111000 : begin
        _zz__zz_regVec_0 = regVec_2168;
      end
      12'b100001111001 : begin
        _zz__zz_regVec_0 = regVec_2169;
      end
      12'b100001111010 : begin
        _zz__zz_regVec_0 = regVec_2170;
      end
      12'b100001111011 : begin
        _zz__zz_regVec_0 = regVec_2171;
      end
      12'b100001111100 : begin
        _zz__zz_regVec_0 = regVec_2172;
      end
      12'b100001111101 : begin
        _zz__zz_regVec_0 = regVec_2173;
      end
      12'b100001111110 : begin
        _zz__zz_regVec_0 = regVec_2174;
      end
      12'b100001111111 : begin
        _zz__zz_regVec_0 = regVec_2175;
      end
      12'b100010000000 : begin
        _zz__zz_regVec_0 = regVec_2176;
      end
      12'b100010000001 : begin
        _zz__zz_regVec_0 = regVec_2177;
      end
      12'b100010000010 : begin
        _zz__zz_regVec_0 = regVec_2178;
      end
      12'b100010000011 : begin
        _zz__zz_regVec_0 = regVec_2179;
      end
      12'b100010000100 : begin
        _zz__zz_regVec_0 = regVec_2180;
      end
      12'b100010000101 : begin
        _zz__zz_regVec_0 = regVec_2181;
      end
      12'b100010000110 : begin
        _zz__zz_regVec_0 = regVec_2182;
      end
      12'b100010000111 : begin
        _zz__zz_regVec_0 = regVec_2183;
      end
      12'b100010001000 : begin
        _zz__zz_regVec_0 = regVec_2184;
      end
      12'b100010001001 : begin
        _zz__zz_regVec_0 = regVec_2185;
      end
      12'b100010001010 : begin
        _zz__zz_regVec_0 = regVec_2186;
      end
      12'b100010001011 : begin
        _zz__zz_regVec_0 = regVec_2187;
      end
      12'b100010001100 : begin
        _zz__zz_regVec_0 = regVec_2188;
      end
      12'b100010001101 : begin
        _zz__zz_regVec_0 = regVec_2189;
      end
      12'b100010001110 : begin
        _zz__zz_regVec_0 = regVec_2190;
      end
      12'b100010001111 : begin
        _zz__zz_regVec_0 = regVec_2191;
      end
      12'b100010010000 : begin
        _zz__zz_regVec_0 = regVec_2192;
      end
      12'b100010010001 : begin
        _zz__zz_regVec_0 = regVec_2193;
      end
      12'b100010010010 : begin
        _zz__zz_regVec_0 = regVec_2194;
      end
      12'b100010010011 : begin
        _zz__zz_regVec_0 = regVec_2195;
      end
      12'b100010010100 : begin
        _zz__zz_regVec_0 = regVec_2196;
      end
      12'b100010010101 : begin
        _zz__zz_regVec_0 = regVec_2197;
      end
      12'b100010010110 : begin
        _zz__zz_regVec_0 = regVec_2198;
      end
      12'b100010010111 : begin
        _zz__zz_regVec_0 = regVec_2199;
      end
      12'b100010011000 : begin
        _zz__zz_regVec_0 = regVec_2200;
      end
      12'b100010011001 : begin
        _zz__zz_regVec_0 = regVec_2201;
      end
      12'b100010011010 : begin
        _zz__zz_regVec_0 = regVec_2202;
      end
      12'b100010011011 : begin
        _zz__zz_regVec_0 = regVec_2203;
      end
      12'b100010011100 : begin
        _zz__zz_regVec_0 = regVec_2204;
      end
      12'b100010011101 : begin
        _zz__zz_regVec_0 = regVec_2205;
      end
      12'b100010011110 : begin
        _zz__zz_regVec_0 = regVec_2206;
      end
      12'b100010011111 : begin
        _zz__zz_regVec_0 = regVec_2207;
      end
      12'b100010100000 : begin
        _zz__zz_regVec_0 = regVec_2208;
      end
      12'b100010100001 : begin
        _zz__zz_regVec_0 = regVec_2209;
      end
      12'b100010100010 : begin
        _zz__zz_regVec_0 = regVec_2210;
      end
      12'b100010100011 : begin
        _zz__zz_regVec_0 = regVec_2211;
      end
      12'b100010100100 : begin
        _zz__zz_regVec_0 = regVec_2212;
      end
      12'b100010100101 : begin
        _zz__zz_regVec_0 = regVec_2213;
      end
      12'b100010100110 : begin
        _zz__zz_regVec_0 = regVec_2214;
      end
      12'b100010100111 : begin
        _zz__zz_regVec_0 = regVec_2215;
      end
      12'b100010101000 : begin
        _zz__zz_regVec_0 = regVec_2216;
      end
      12'b100010101001 : begin
        _zz__zz_regVec_0 = regVec_2217;
      end
      12'b100010101010 : begin
        _zz__zz_regVec_0 = regVec_2218;
      end
      12'b100010101011 : begin
        _zz__zz_regVec_0 = regVec_2219;
      end
      12'b100010101100 : begin
        _zz__zz_regVec_0 = regVec_2220;
      end
      12'b100010101101 : begin
        _zz__zz_regVec_0 = regVec_2221;
      end
      12'b100010101110 : begin
        _zz__zz_regVec_0 = regVec_2222;
      end
      12'b100010101111 : begin
        _zz__zz_regVec_0 = regVec_2223;
      end
      12'b100010110000 : begin
        _zz__zz_regVec_0 = regVec_2224;
      end
      12'b100010110001 : begin
        _zz__zz_regVec_0 = regVec_2225;
      end
      12'b100010110010 : begin
        _zz__zz_regVec_0 = regVec_2226;
      end
      12'b100010110011 : begin
        _zz__zz_regVec_0 = regVec_2227;
      end
      12'b100010110100 : begin
        _zz__zz_regVec_0 = regVec_2228;
      end
      12'b100010110101 : begin
        _zz__zz_regVec_0 = regVec_2229;
      end
      12'b100010110110 : begin
        _zz__zz_regVec_0 = regVec_2230;
      end
      12'b100010110111 : begin
        _zz__zz_regVec_0 = regVec_2231;
      end
      12'b100010111000 : begin
        _zz__zz_regVec_0 = regVec_2232;
      end
      12'b100010111001 : begin
        _zz__zz_regVec_0 = regVec_2233;
      end
      12'b100010111010 : begin
        _zz__zz_regVec_0 = regVec_2234;
      end
      12'b100010111011 : begin
        _zz__zz_regVec_0 = regVec_2235;
      end
      12'b100010111100 : begin
        _zz__zz_regVec_0 = regVec_2236;
      end
      12'b100010111101 : begin
        _zz__zz_regVec_0 = regVec_2237;
      end
      12'b100010111110 : begin
        _zz__zz_regVec_0 = regVec_2238;
      end
      12'b100010111111 : begin
        _zz__zz_regVec_0 = regVec_2239;
      end
      12'b100011000000 : begin
        _zz__zz_regVec_0 = regVec_2240;
      end
      12'b100011000001 : begin
        _zz__zz_regVec_0 = regVec_2241;
      end
      12'b100011000010 : begin
        _zz__zz_regVec_0 = regVec_2242;
      end
      12'b100011000011 : begin
        _zz__zz_regVec_0 = regVec_2243;
      end
      12'b100011000100 : begin
        _zz__zz_regVec_0 = regVec_2244;
      end
      12'b100011000101 : begin
        _zz__zz_regVec_0 = regVec_2245;
      end
      12'b100011000110 : begin
        _zz__zz_regVec_0 = regVec_2246;
      end
      12'b100011000111 : begin
        _zz__zz_regVec_0 = regVec_2247;
      end
      12'b100011001000 : begin
        _zz__zz_regVec_0 = regVec_2248;
      end
      12'b100011001001 : begin
        _zz__zz_regVec_0 = regVec_2249;
      end
      12'b100011001010 : begin
        _zz__zz_regVec_0 = regVec_2250;
      end
      12'b100011001011 : begin
        _zz__zz_regVec_0 = regVec_2251;
      end
      12'b100011001100 : begin
        _zz__zz_regVec_0 = regVec_2252;
      end
      12'b100011001101 : begin
        _zz__zz_regVec_0 = regVec_2253;
      end
      12'b100011001110 : begin
        _zz__zz_regVec_0 = regVec_2254;
      end
      12'b100011001111 : begin
        _zz__zz_regVec_0 = regVec_2255;
      end
      12'b100011010000 : begin
        _zz__zz_regVec_0 = regVec_2256;
      end
      12'b100011010001 : begin
        _zz__zz_regVec_0 = regVec_2257;
      end
      12'b100011010010 : begin
        _zz__zz_regVec_0 = regVec_2258;
      end
      12'b100011010011 : begin
        _zz__zz_regVec_0 = regVec_2259;
      end
      12'b100011010100 : begin
        _zz__zz_regVec_0 = regVec_2260;
      end
      12'b100011010101 : begin
        _zz__zz_regVec_0 = regVec_2261;
      end
      12'b100011010110 : begin
        _zz__zz_regVec_0 = regVec_2262;
      end
      12'b100011010111 : begin
        _zz__zz_regVec_0 = regVec_2263;
      end
      12'b100011011000 : begin
        _zz__zz_regVec_0 = regVec_2264;
      end
      12'b100011011001 : begin
        _zz__zz_regVec_0 = regVec_2265;
      end
      12'b100011011010 : begin
        _zz__zz_regVec_0 = regVec_2266;
      end
      12'b100011011011 : begin
        _zz__zz_regVec_0 = regVec_2267;
      end
      12'b100011011100 : begin
        _zz__zz_regVec_0 = regVec_2268;
      end
      12'b100011011101 : begin
        _zz__zz_regVec_0 = regVec_2269;
      end
      12'b100011011110 : begin
        _zz__zz_regVec_0 = regVec_2270;
      end
      12'b100011011111 : begin
        _zz__zz_regVec_0 = regVec_2271;
      end
      12'b100011100000 : begin
        _zz__zz_regVec_0 = regVec_2272;
      end
      12'b100011100001 : begin
        _zz__zz_regVec_0 = regVec_2273;
      end
      12'b100011100010 : begin
        _zz__zz_regVec_0 = regVec_2274;
      end
      12'b100011100011 : begin
        _zz__zz_regVec_0 = regVec_2275;
      end
      12'b100011100100 : begin
        _zz__zz_regVec_0 = regVec_2276;
      end
      12'b100011100101 : begin
        _zz__zz_regVec_0 = regVec_2277;
      end
      12'b100011100110 : begin
        _zz__zz_regVec_0 = regVec_2278;
      end
      12'b100011100111 : begin
        _zz__zz_regVec_0 = regVec_2279;
      end
      12'b100011101000 : begin
        _zz__zz_regVec_0 = regVec_2280;
      end
      12'b100011101001 : begin
        _zz__zz_regVec_0 = regVec_2281;
      end
      12'b100011101010 : begin
        _zz__zz_regVec_0 = regVec_2282;
      end
      12'b100011101011 : begin
        _zz__zz_regVec_0 = regVec_2283;
      end
      12'b100011101100 : begin
        _zz__zz_regVec_0 = regVec_2284;
      end
      12'b100011101101 : begin
        _zz__zz_regVec_0 = regVec_2285;
      end
      12'b100011101110 : begin
        _zz__zz_regVec_0 = regVec_2286;
      end
      12'b100011101111 : begin
        _zz__zz_regVec_0 = regVec_2287;
      end
      12'b100011110000 : begin
        _zz__zz_regVec_0 = regVec_2288;
      end
      12'b100011110001 : begin
        _zz__zz_regVec_0 = regVec_2289;
      end
      12'b100011110010 : begin
        _zz__zz_regVec_0 = regVec_2290;
      end
      12'b100011110011 : begin
        _zz__zz_regVec_0 = regVec_2291;
      end
      12'b100011110100 : begin
        _zz__zz_regVec_0 = regVec_2292;
      end
      12'b100011110101 : begin
        _zz__zz_regVec_0 = regVec_2293;
      end
      12'b100011110110 : begin
        _zz__zz_regVec_0 = regVec_2294;
      end
      12'b100011110111 : begin
        _zz__zz_regVec_0 = regVec_2295;
      end
      12'b100011111000 : begin
        _zz__zz_regVec_0 = regVec_2296;
      end
      12'b100011111001 : begin
        _zz__zz_regVec_0 = regVec_2297;
      end
      12'b100011111010 : begin
        _zz__zz_regVec_0 = regVec_2298;
      end
      12'b100011111011 : begin
        _zz__zz_regVec_0 = regVec_2299;
      end
      12'b100011111100 : begin
        _zz__zz_regVec_0 = regVec_2300;
      end
      12'b100011111101 : begin
        _zz__zz_regVec_0 = regVec_2301;
      end
      12'b100011111110 : begin
        _zz__zz_regVec_0 = regVec_2302;
      end
      12'b100011111111 : begin
        _zz__zz_regVec_0 = regVec_2303;
      end
      12'b100100000000 : begin
        _zz__zz_regVec_0 = regVec_2304;
      end
      12'b100100000001 : begin
        _zz__zz_regVec_0 = regVec_2305;
      end
      12'b100100000010 : begin
        _zz__zz_regVec_0 = regVec_2306;
      end
      12'b100100000011 : begin
        _zz__zz_regVec_0 = regVec_2307;
      end
      12'b100100000100 : begin
        _zz__zz_regVec_0 = regVec_2308;
      end
      12'b100100000101 : begin
        _zz__zz_regVec_0 = regVec_2309;
      end
      12'b100100000110 : begin
        _zz__zz_regVec_0 = regVec_2310;
      end
      12'b100100000111 : begin
        _zz__zz_regVec_0 = regVec_2311;
      end
      12'b100100001000 : begin
        _zz__zz_regVec_0 = regVec_2312;
      end
      12'b100100001001 : begin
        _zz__zz_regVec_0 = regVec_2313;
      end
      12'b100100001010 : begin
        _zz__zz_regVec_0 = regVec_2314;
      end
      12'b100100001011 : begin
        _zz__zz_regVec_0 = regVec_2315;
      end
      12'b100100001100 : begin
        _zz__zz_regVec_0 = regVec_2316;
      end
      12'b100100001101 : begin
        _zz__zz_regVec_0 = regVec_2317;
      end
      12'b100100001110 : begin
        _zz__zz_regVec_0 = regVec_2318;
      end
      12'b100100001111 : begin
        _zz__zz_regVec_0 = regVec_2319;
      end
      12'b100100010000 : begin
        _zz__zz_regVec_0 = regVec_2320;
      end
      12'b100100010001 : begin
        _zz__zz_regVec_0 = regVec_2321;
      end
      12'b100100010010 : begin
        _zz__zz_regVec_0 = regVec_2322;
      end
      12'b100100010011 : begin
        _zz__zz_regVec_0 = regVec_2323;
      end
      12'b100100010100 : begin
        _zz__zz_regVec_0 = regVec_2324;
      end
      12'b100100010101 : begin
        _zz__zz_regVec_0 = regVec_2325;
      end
      12'b100100010110 : begin
        _zz__zz_regVec_0 = regVec_2326;
      end
      12'b100100010111 : begin
        _zz__zz_regVec_0 = regVec_2327;
      end
      12'b100100011000 : begin
        _zz__zz_regVec_0 = regVec_2328;
      end
      12'b100100011001 : begin
        _zz__zz_regVec_0 = regVec_2329;
      end
      12'b100100011010 : begin
        _zz__zz_regVec_0 = regVec_2330;
      end
      12'b100100011011 : begin
        _zz__zz_regVec_0 = regVec_2331;
      end
      12'b100100011100 : begin
        _zz__zz_regVec_0 = regVec_2332;
      end
      12'b100100011101 : begin
        _zz__zz_regVec_0 = regVec_2333;
      end
      12'b100100011110 : begin
        _zz__zz_regVec_0 = regVec_2334;
      end
      12'b100100011111 : begin
        _zz__zz_regVec_0 = regVec_2335;
      end
      12'b100100100000 : begin
        _zz__zz_regVec_0 = regVec_2336;
      end
      12'b100100100001 : begin
        _zz__zz_regVec_0 = regVec_2337;
      end
      12'b100100100010 : begin
        _zz__zz_regVec_0 = regVec_2338;
      end
      12'b100100100011 : begin
        _zz__zz_regVec_0 = regVec_2339;
      end
      12'b100100100100 : begin
        _zz__zz_regVec_0 = regVec_2340;
      end
      12'b100100100101 : begin
        _zz__zz_regVec_0 = regVec_2341;
      end
      12'b100100100110 : begin
        _zz__zz_regVec_0 = regVec_2342;
      end
      12'b100100100111 : begin
        _zz__zz_regVec_0 = regVec_2343;
      end
      12'b100100101000 : begin
        _zz__zz_regVec_0 = regVec_2344;
      end
      12'b100100101001 : begin
        _zz__zz_regVec_0 = regVec_2345;
      end
      12'b100100101010 : begin
        _zz__zz_regVec_0 = regVec_2346;
      end
      12'b100100101011 : begin
        _zz__zz_regVec_0 = regVec_2347;
      end
      12'b100100101100 : begin
        _zz__zz_regVec_0 = regVec_2348;
      end
      12'b100100101101 : begin
        _zz__zz_regVec_0 = regVec_2349;
      end
      12'b100100101110 : begin
        _zz__zz_regVec_0 = regVec_2350;
      end
      12'b100100101111 : begin
        _zz__zz_regVec_0 = regVec_2351;
      end
      12'b100100110000 : begin
        _zz__zz_regVec_0 = regVec_2352;
      end
      12'b100100110001 : begin
        _zz__zz_regVec_0 = regVec_2353;
      end
      12'b100100110010 : begin
        _zz__zz_regVec_0 = regVec_2354;
      end
      12'b100100110011 : begin
        _zz__zz_regVec_0 = regVec_2355;
      end
      12'b100100110100 : begin
        _zz__zz_regVec_0 = regVec_2356;
      end
      12'b100100110101 : begin
        _zz__zz_regVec_0 = regVec_2357;
      end
      12'b100100110110 : begin
        _zz__zz_regVec_0 = regVec_2358;
      end
      12'b100100110111 : begin
        _zz__zz_regVec_0 = regVec_2359;
      end
      12'b100100111000 : begin
        _zz__zz_regVec_0 = regVec_2360;
      end
      12'b100100111001 : begin
        _zz__zz_regVec_0 = regVec_2361;
      end
      12'b100100111010 : begin
        _zz__zz_regVec_0 = regVec_2362;
      end
      12'b100100111011 : begin
        _zz__zz_regVec_0 = regVec_2363;
      end
      12'b100100111100 : begin
        _zz__zz_regVec_0 = regVec_2364;
      end
      12'b100100111101 : begin
        _zz__zz_regVec_0 = regVec_2365;
      end
      12'b100100111110 : begin
        _zz__zz_regVec_0 = regVec_2366;
      end
      12'b100100111111 : begin
        _zz__zz_regVec_0 = regVec_2367;
      end
      12'b100101000000 : begin
        _zz__zz_regVec_0 = regVec_2368;
      end
      12'b100101000001 : begin
        _zz__zz_regVec_0 = regVec_2369;
      end
      12'b100101000010 : begin
        _zz__zz_regVec_0 = regVec_2370;
      end
      12'b100101000011 : begin
        _zz__zz_regVec_0 = regVec_2371;
      end
      12'b100101000100 : begin
        _zz__zz_regVec_0 = regVec_2372;
      end
      12'b100101000101 : begin
        _zz__zz_regVec_0 = regVec_2373;
      end
      12'b100101000110 : begin
        _zz__zz_regVec_0 = regVec_2374;
      end
      12'b100101000111 : begin
        _zz__zz_regVec_0 = regVec_2375;
      end
      12'b100101001000 : begin
        _zz__zz_regVec_0 = regVec_2376;
      end
      12'b100101001001 : begin
        _zz__zz_regVec_0 = regVec_2377;
      end
      12'b100101001010 : begin
        _zz__zz_regVec_0 = regVec_2378;
      end
      12'b100101001011 : begin
        _zz__zz_regVec_0 = regVec_2379;
      end
      12'b100101001100 : begin
        _zz__zz_regVec_0 = regVec_2380;
      end
      12'b100101001101 : begin
        _zz__zz_regVec_0 = regVec_2381;
      end
      12'b100101001110 : begin
        _zz__zz_regVec_0 = regVec_2382;
      end
      12'b100101001111 : begin
        _zz__zz_regVec_0 = regVec_2383;
      end
      12'b100101010000 : begin
        _zz__zz_regVec_0 = regVec_2384;
      end
      12'b100101010001 : begin
        _zz__zz_regVec_0 = regVec_2385;
      end
      12'b100101010010 : begin
        _zz__zz_regVec_0 = regVec_2386;
      end
      12'b100101010011 : begin
        _zz__zz_regVec_0 = regVec_2387;
      end
      12'b100101010100 : begin
        _zz__zz_regVec_0 = regVec_2388;
      end
      12'b100101010101 : begin
        _zz__zz_regVec_0 = regVec_2389;
      end
      12'b100101010110 : begin
        _zz__zz_regVec_0 = regVec_2390;
      end
      12'b100101010111 : begin
        _zz__zz_regVec_0 = regVec_2391;
      end
      12'b100101011000 : begin
        _zz__zz_regVec_0 = regVec_2392;
      end
      12'b100101011001 : begin
        _zz__zz_regVec_0 = regVec_2393;
      end
      12'b100101011010 : begin
        _zz__zz_regVec_0 = regVec_2394;
      end
      12'b100101011011 : begin
        _zz__zz_regVec_0 = regVec_2395;
      end
      12'b100101011100 : begin
        _zz__zz_regVec_0 = regVec_2396;
      end
      12'b100101011101 : begin
        _zz__zz_regVec_0 = regVec_2397;
      end
      12'b100101011110 : begin
        _zz__zz_regVec_0 = regVec_2398;
      end
      12'b100101011111 : begin
        _zz__zz_regVec_0 = regVec_2399;
      end
      12'b100101100000 : begin
        _zz__zz_regVec_0 = regVec_2400;
      end
      12'b100101100001 : begin
        _zz__zz_regVec_0 = regVec_2401;
      end
      12'b100101100010 : begin
        _zz__zz_regVec_0 = regVec_2402;
      end
      12'b100101100011 : begin
        _zz__zz_regVec_0 = regVec_2403;
      end
      12'b100101100100 : begin
        _zz__zz_regVec_0 = regVec_2404;
      end
      12'b100101100101 : begin
        _zz__zz_regVec_0 = regVec_2405;
      end
      12'b100101100110 : begin
        _zz__zz_regVec_0 = regVec_2406;
      end
      12'b100101100111 : begin
        _zz__zz_regVec_0 = regVec_2407;
      end
      12'b100101101000 : begin
        _zz__zz_regVec_0 = regVec_2408;
      end
      12'b100101101001 : begin
        _zz__zz_regVec_0 = regVec_2409;
      end
      12'b100101101010 : begin
        _zz__zz_regVec_0 = regVec_2410;
      end
      12'b100101101011 : begin
        _zz__zz_regVec_0 = regVec_2411;
      end
      12'b100101101100 : begin
        _zz__zz_regVec_0 = regVec_2412;
      end
      12'b100101101101 : begin
        _zz__zz_regVec_0 = regVec_2413;
      end
      12'b100101101110 : begin
        _zz__zz_regVec_0 = regVec_2414;
      end
      12'b100101101111 : begin
        _zz__zz_regVec_0 = regVec_2415;
      end
      12'b100101110000 : begin
        _zz__zz_regVec_0 = regVec_2416;
      end
      12'b100101110001 : begin
        _zz__zz_regVec_0 = regVec_2417;
      end
      12'b100101110010 : begin
        _zz__zz_regVec_0 = regVec_2418;
      end
      12'b100101110011 : begin
        _zz__zz_regVec_0 = regVec_2419;
      end
      12'b100101110100 : begin
        _zz__zz_regVec_0 = regVec_2420;
      end
      12'b100101110101 : begin
        _zz__zz_regVec_0 = regVec_2421;
      end
      12'b100101110110 : begin
        _zz__zz_regVec_0 = regVec_2422;
      end
      12'b100101110111 : begin
        _zz__zz_regVec_0 = regVec_2423;
      end
      12'b100101111000 : begin
        _zz__zz_regVec_0 = regVec_2424;
      end
      12'b100101111001 : begin
        _zz__zz_regVec_0 = regVec_2425;
      end
      12'b100101111010 : begin
        _zz__zz_regVec_0 = regVec_2426;
      end
      12'b100101111011 : begin
        _zz__zz_regVec_0 = regVec_2427;
      end
      12'b100101111100 : begin
        _zz__zz_regVec_0 = regVec_2428;
      end
      12'b100101111101 : begin
        _zz__zz_regVec_0 = regVec_2429;
      end
      12'b100101111110 : begin
        _zz__zz_regVec_0 = regVec_2430;
      end
      12'b100101111111 : begin
        _zz__zz_regVec_0 = regVec_2431;
      end
      12'b100110000000 : begin
        _zz__zz_regVec_0 = regVec_2432;
      end
      12'b100110000001 : begin
        _zz__zz_regVec_0 = regVec_2433;
      end
      12'b100110000010 : begin
        _zz__zz_regVec_0 = regVec_2434;
      end
      12'b100110000011 : begin
        _zz__zz_regVec_0 = regVec_2435;
      end
      12'b100110000100 : begin
        _zz__zz_regVec_0 = regVec_2436;
      end
      12'b100110000101 : begin
        _zz__zz_regVec_0 = regVec_2437;
      end
      12'b100110000110 : begin
        _zz__zz_regVec_0 = regVec_2438;
      end
      12'b100110000111 : begin
        _zz__zz_regVec_0 = regVec_2439;
      end
      12'b100110001000 : begin
        _zz__zz_regVec_0 = regVec_2440;
      end
      12'b100110001001 : begin
        _zz__zz_regVec_0 = regVec_2441;
      end
      12'b100110001010 : begin
        _zz__zz_regVec_0 = regVec_2442;
      end
      12'b100110001011 : begin
        _zz__zz_regVec_0 = regVec_2443;
      end
      12'b100110001100 : begin
        _zz__zz_regVec_0 = regVec_2444;
      end
      12'b100110001101 : begin
        _zz__zz_regVec_0 = regVec_2445;
      end
      12'b100110001110 : begin
        _zz__zz_regVec_0 = regVec_2446;
      end
      12'b100110001111 : begin
        _zz__zz_regVec_0 = regVec_2447;
      end
      12'b100110010000 : begin
        _zz__zz_regVec_0 = regVec_2448;
      end
      12'b100110010001 : begin
        _zz__zz_regVec_0 = regVec_2449;
      end
      12'b100110010010 : begin
        _zz__zz_regVec_0 = regVec_2450;
      end
      12'b100110010011 : begin
        _zz__zz_regVec_0 = regVec_2451;
      end
      12'b100110010100 : begin
        _zz__zz_regVec_0 = regVec_2452;
      end
      12'b100110010101 : begin
        _zz__zz_regVec_0 = regVec_2453;
      end
      12'b100110010110 : begin
        _zz__zz_regVec_0 = regVec_2454;
      end
      12'b100110010111 : begin
        _zz__zz_regVec_0 = regVec_2455;
      end
      12'b100110011000 : begin
        _zz__zz_regVec_0 = regVec_2456;
      end
      12'b100110011001 : begin
        _zz__zz_regVec_0 = regVec_2457;
      end
      12'b100110011010 : begin
        _zz__zz_regVec_0 = regVec_2458;
      end
      12'b100110011011 : begin
        _zz__zz_regVec_0 = regVec_2459;
      end
      12'b100110011100 : begin
        _zz__zz_regVec_0 = regVec_2460;
      end
      12'b100110011101 : begin
        _zz__zz_regVec_0 = regVec_2461;
      end
      12'b100110011110 : begin
        _zz__zz_regVec_0 = regVec_2462;
      end
      12'b100110011111 : begin
        _zz__zz_regVec_0 = regVec_2463;
      end
      12'b100110100000 : begin
        _zz__zz_regVec_0 = regVec_2464;
      end
      12'b100110100001 : begin
        _zz__zz_regVec_0 = regVec_2465;
      end
      12'b100110100010 : begin
        _zz__zz_regVec_0 = regVec_2466;
      end
      12'b100110100011 : begin
        _zz__zz_regVec_0 = regVec_2467;
      end
      12'b100110100100 : begin
        _zz__zz_regVec_0 = regVec_2468;
      end
      12'b100110100101 : begin
        _zz__zz_regVec_0 = regVec_2469;
      end
      12'b100110100110 : begin
        _zz__zz_regVec_0 = regVec_2470;
      end
      12'b100110100111 : begin
        _zz__zz_regVec_0 = regVec_2471;
      end
      12'b100110101000 : begin
        _zz__zz_regVec_0 = regVec_2472;
      end
      12'b100110101001 : begin
        _zz__zz_regVec_0 = regVec_2473;
      end
      12'b100110101010 : begin
        _zz__zz_regVec_0 = regVec_2474;
      end
      12'b100110101011 : begin
        _zz__zz_regVec_0 = regVec_2475;
      end
      12'b100110101100 : begin
        _zz__zz_regVec_0 = regVec_2476;
      end
      12'b100110101101 : begin
        _zz__zz_regVec_0 = regVec_2477;
      end
      12'b100110101110 : begin
        _zz__zz_regVec_0 = regVec_2478;
      end
      12'b100110101111 : begin
        _zz__zz_regVec_0 = regVec_2479;
      end
      12'b100110110000 : begin
        _zz__zz_regVec_0 = regVec_2480;
      end
      12'b100110110001 : begin
        _zz__zz_regVec_0 = regVec_2481;
      end
      12'b100110110010 : begin
        _zz__zz_regVec_0 = regVec_2482;
      end
      12'b100110110011 : begin
        _zz__zz_regVec_0 = regVec_2483;
      end
      12'b100110110100 : begin
        _zz__zz_regVec_0 = regVec_2484;
      end
      12'b100110110101 : begin
        _zz__zz_regVec_0 = regVec_2485;
      end
      12'b100110110110 : begin
        _zz__zz_regVec_0 = regVec_2486;
      end
      12'b100110110111 : begin
        _zz__zz_regVec_0 = regVec_2487;
      end
      12'b100110111000 : begin
        _zz__zz_regVec_0 = regVec_2488;
      end
      12'b100110111001 : begin
        _zz__zz_regVec_0 = regVec_2489;
      end
      12'b100110111010 : begin
        _zz__zz_regVec_0 = regVec_2490;
      end
      12'b100110111011 : begin
        _zz__zz_regVec_0 = regVec_2491;
      end
      12'b100110111100 : begin
        _zz__zz_regVec_0 = regVec_2492;
      end
      12'b100110111101 : begin
        _zz__zz_regVec_0 = regVec_2493;
      end
      12'b100110111110 : begin
        _zz__zz_regVec_0 = regVec_2494;
      end
      12'b100110111111 : begin
        _zz__zz_regVec_0 = regVec_2495;
      end
      12'b100111000000 : begin
        _zz__zz_regVec_0 = regVec_2496;
      end
      12'b100111000001 : begin
        _zz__zz_regVec_0 = regVec_2497;
      end
      12'b100111000010 : begin
        _zz__zz_regVec_0 = regVec_2498;
      end
      12'b100111000011 : begin
        _zz__zz_regVec_0 = regVec_2499;
      end
      12'b100111000100 : begin
        _zz__zz_regVec_0 = regVec_2500;
      end
      12'b100111000101 : begin
        _zz__zz_regVec_0 = regVec_2501;
      end
      12'b100111000110 : begin
        _zz__zz_regVec_0 = regVec_2502;
      end
      12'b100111000111 : begin
        _zz__zz_regVec_0 = regVec_2503;
      end
      12'b100111001000 : begin
        _zz__zz_regVec_0 = regVec_2504;
      end
      12'b100111001001 : begin
        _zz__zz_regVec_0 = regVec_2505;
      end
      12'b100111001010 : begin
        _zz__zz_regVec_0 = regVec_2506;
      end
      12'b100111001011 : begin
        _zz__zz_regVec_0 = regVec_2507;
      end
      12'b100111001100 : begin
        _zz__zz_regVec_0 = regVec_2508;
      end
      12'b100111001101 : begin
        _zz__zz_regVec_0 = regVec_2509;
      end
      12'b100111001110 : begin
        _zz__zz_regVec_0 = regVec_2510;
      end
      12'b100111001111 : begin
        _zz__zz_regVec_0 = regVec_2511;
      end
      12'b100111010000 : begin
        _zz__zz_regVec_0 = regVec_2512;
      end
      12'b100111010001 : begin
        _zz__zz_regVec_0 = regVec_2513;
      end
      12'b100111010010 : begin
        _zz__zz_regVec_0 = regVec_2514;
      end
      12'b100111010011 : begin
        _zz__zz_regVec_0 = regVec_2515;
      end
      12'b100111010100 : begin
        _zz__zz_regVec_0 = regVec_2516;
      end
      12'b100111010101 : begin
        _zz__zz_regVec_0 = regVec_2517;
      end
      12'b100111010110 : begin
        _zz__zz_regVec_0 = regVec_2518;
      end
      12'b100111010111 : begin
        _zz__zz_regVec_0 = regVec_2519;
      end
      12'b100111011000 : begin
        _zz__zz_regVec_0 = regVec_2520;
      end
      12'b100111011001 : begin
        _zz__zz_regVec_0 = regVec_2521;
      end
      12'b100111011010 : begin
        _zz__zz_regVec_0 = regVec_2522;
      end
      12'b100111011011 : begin
        _zz__zz_regVec_0 = regVec_2523;
      end
      12'b100111011100 : begin
        _zz__zz_regVec_0 = regVec_2524;
      end
      12'b100111011101 : begin
        _zz__zz_regVec_0 = regVec_2525;
      end
      12'b100111011110 : begin
        _zz__zz_regVec_0 = regVec_2526;
      end
      12'b100111011111 : begin
        _zz__zz_regVec_0 = regVec_2527;
      end
      12'b100111100000 : begin
        _zz__zz_regVec_0 = regVec_2528;
      end
      12'b100111100001 : begin
        _zz__zz_regVec_0 = regVec_2529;
      end
      12'b100111100010 : begin
        _zz__zz_regVec_0 = regVec_2530;
      end
      12'b100111100011 : begin
        _zz__zz_regVec_0 = regVec_2531;
      end
      12'b100111100100 : begin
        _zz__zz_regVec_0 = regVec_2532;
      end
      12'b100111100101 : begin
        _zz__zz_regVec_0 = regVec_2533;
      end
      12'b100111100110 : begin
        _zz__zz_regVec_0 = regVec_2534;
      end
      12'b100111100111 : begin
        _zz__zz_regVec_0 = regVec_2535;
      end
      12'b100111101000 : begin
        _zz__zz_regVec_0 = regVec_2536;
      end
      12'b100111101001 : begin
        _zz__zz_regVec_0 = regVec_2537;
      end
      12'b100111101010 : begin
        _zz__zz_regVec_0 = regVec_2538;
      end
      12'b100111101011 : begin
        _zz__zz_regVec_0 = regVec_2539;
      end
      12'b100111101100 : begin
        _zz__zz_regVec_0 = regVec_2540;
      end
      12'b100111101101 : begin
        _zz__zz_regVec_0 = regVec_2541;
      end
      12'b100111101110 : begin
        _zz__zz_regVec_0 = regVec_2542;
      end
      12'b100111101111 : begin
        _zz__zz_regVec_0 = regVec_2543;
      end
      12'b100111110000 : begin
        _zz__zz_regVec_0 = regVec_2544;
      end
      12'b100111110001 : begin
        _zz__zz_regVec_0 = regVec_2545;
      end
      12'b100111110010 : begin
        _zz__zz_regVec_0 = regVec_2546;
      end
      12'b100111110011 : begin
        _zz__zz_regVec_0 = regVec_2547;
      end
      12'b100111110100 : begin
        _zz__zz_regVec_0 = regVec_2548;
      end
      12'b100111110101 : begin
        _zz__zz_regVec_0 = regVec_2549;
      end
      12'b100111110110 : begin
        _zz__zz_regVec_0 = regVec_2550;
      end
      12'b100111110111 : begin
        _zz__zz_regVec_0 = regVec_2551;
      end
      12'b100111111000 : begin
        _zz__zz_regVec_0 = regVec_2552;
      end
      12'b100111111001 : begin
        _zz__zz_regVec_0 = regVec_2553;
      end
      12'b100111111010 : begin
        _zz__zz_regVec_0 = regVec_2554;
      end
      12'b100111111011 : begin
        _zz__zz_regVec_0 = regVec_2555;
      end
      12'b100111111100 : begin
        _zz__zz_regVec_0 = regVec_2556;
      end
      12'b100111111101 : begin
        _zz__zz_regVec_0 = regVec_2557;
      end
      12'b100111111110 : begin
        _zz__zz_regVec_0 = regVec_2558;
      end
      12'b100111111111 : begin
        _zz__zz_regVec_0 = regVec_2559;
      end
      12'b101000000000 : begin
        _zz__zz_regVec_0 = regVec_2560;
      end
      12'b101000000001 : begin
        _zz__zz_regVec_0 = regVec_2561;
      end
      12'b101000000010 : begin
        _zz__zz_regVec_0 = regVec_2562;
      end
      12'b101000000011 : begin
        _zz__zz_regVec_0 = regVec_2563;
      end
      12'b101000000100 : begin
        _zz__zz_regVec_0 = regVec_2564;
      end
      12'b101000000101 : begin
        _zz__zz_regVec_0 = regVec_2565;
      end
      12'b101000000110 : begin
        _zz__zz_regVec_0 = regVec_2566;
      end
      12'b101000000111 : begin
        _zz__zz_regVec_0 = regVec_2567;
      end
      12'b101000001000 : begin
        _zz__zz_regVec_0 = regVec_2568;
      end
      12'b101000001001 : begin
        _zz__zz_regVec_0 = regVec_2569;
      end
      12'b101000001010 : begin
        _zz__zz_regVec_0 = regVec_2570;
      end
      12'b101000001011 : begin
        _zz__zz_regVec_0 = regVec_2571;
      end
      12'b101000001100 : begin
        _zz__zz_regVec_0 = regVec_2572;
      end
      12'b101000001101 : begin
        _zz__zz_regVec_0 = regVec_2573;
      end
      12'b101000001110 : begin
        _zz__zz_regVec_0 = regVec_2574;
      end
      12'b101000001111 : begin
        _zz__zz_regVec_0 = regVec_2575;
      end
      12'b101000010000 : begin
        _zz__zz_regVec_0 = regVec_2576;
      end
      12'b101000010001 : begin
        _zz__zz_regVec_0 = regVec_2577;
      end
      12'b101000010010 : begin
        _zz__zz_regVec_0 = regVec_2578;
      end
      12'b101000010011 : begin
        _zz__zz_regVec_0 = regVec_2579;
      end
      12'b101000010100 : begin
        _zz__zz_regVec_0 = regVec_2580;
      end
      12'b101000010101 : begin
        _zz__zz_regVec_0 = regVec_2581;
      end
      12'b101000010110 : begin
        _zz__zz_regVec_0 = regVec_2582;
      end
      12'b101000010111 : begin
        _zz__zz_regVec_0 = regVec_2583;
      end
      12'b101000011000 : begin
        _zz__zz_regVec_0 = regVec_2584;
      end
      12'b101000011001 : begin
        _zz__zz_regVec_0 = regVec_2585;
      end
      12'b101000011010 : begin
        _zz__zz_regVec_0 = regVec_2586;
      end
      12'b101000011011 : begin
        _zz__zz_regVec_0 = regVec_2587;
      end
      12'b101000011100 : begin
        _zz__zz_regVec_0 = regVec_2588;
      end
      12'b101000011101 : begin
        _zz__zz_regVec_0 = regVec_2589;
      end
      12'b101000011110 : begin
        _zz__zz_regVec_0 = regVec_2590;
      end
      12'b101000011111 : begin
        _zz__zz_regVec_0 = regVec_2591;
      end
      12'b101000100000 : begin
        _zz__zz_regVec_0 = regVec_2592;
      end
      12'b101000100001 : begin
        _zz__zz_regVec_0 = regVec_2593;
      end
      12'b101000100010 : begin
        _zz__zz_regVec_0 = regVec_2594;
      end
      12'b101000100011 : begin
        _zz__zz_regVec_0 = regVec_2595;
      end
      12'b101000100100 : begin
        _zz__zz_regVec_0 = regVec_2596;
      end
      12'b101000100101 : begin
        _zz__zz_regVec_0 = regVec_2597;
      end
      12'b101000100110 : begin
        _zz__zz_regVec_0 = regVec_2598;
      end
      12'b101000100111 : begin
        _zz__zz_regVec_0 = regVec_2599;
      end
      12'b101000101000 : begin
        _zz__zz_regVec_0 = regVec_2600;
      end
      12'b101000101001 : begin
        _zz__zz_regVec_0 = regVec_2601;
      end
      12'b101000101010 : begin
        _zz__zz_regVec_0 = regVec_2602;
      end
      12'b101000101011 : begin
        _zz__zz_regVec_0 = regVec_2603;
      end
      12'b101000101100 : begin
        _zz__zz_regVec_0 = regVec_2604;
      end
      12'b101000101101 : begin
        _zz__zz_regVec_0 = regVec_2605;
      end
      12'b101000101110 : begin
        _zz__zz_regVec_0 = regVec_2606;
      end
      12'b101000101111 : begin
        _zz__zz_regVec_0 = regVec_2607;
      end
      12'b101000110000 : begin
        _zz__zz_regVec_0 = regVec_2608;
      end
      12'b101000110001 : begin
        _zz__zz_regVec_0 = regVec_2609;
      end
      12'b101000110010 : begin
        _zz__zz_regVec_0 = regVec_2610;
      end
      12'b101000110011 : begin
        _zz__zz_regVec_0 = regVec_2611;
      end
      12'b101000110100 : begin
        _zz__zz_regVec_0 = regVec_2612;
      end
      12'b101000110101 : begin
        _zz__zz_regVec_0 = regVec_2613;
      end
      12'b101000110110 : begin
        _zz__zz_regVec_0 = regVec_2614;
      end
      12'b101000110111 : begin
        _zz__zz_regVec_0 = regVec_2615;
      end
      12'b101000111000 : begin
        _zz__zz_regVec_0 = regVec_2616;
      end
      12'b101000111001 : begin
        _zz__zz_regVec_0 = regVec_2617;
      end
      12'b101000111010 : begin
        _zz__zz_regVec_0 = regVec_2618;
      end
      12'b101000111011 : begin
        _zz__zz_regVec_0 = regVec_2619;
      end
      12'b101000111100 : begin
        _zz__zz_regVec_0 = regVec_2620;
      end
      12'b101000111101 : begin
        _zz__zz_regVec_0 = regVec_2621;
      end
      12'b101000111110 : begin
        _zz__zz_regVec_0 = regVec_2622;
      end
      12'b101000111111 : begin
        _zz__zz_regVec_0 = regVec_2623;
      end
      12'b101001000000 : begin
        _zz__zz_regVec_0 = regVec_2624;
      end
      12'b101001000001 : begin
        _zz__zz_regVec_0 = regVec_2625;
      end
      12'b101001000010 : begin
        _zz__zz_regVec_0 = regVec_2626;
      end
      12'b101001000011 : begin
        _zz__zz_regVec_0 = regVec_2627;
      end
      12'b101001000100 : begin
        _zz__zz_regVec_0 = regVec_2628;
      end
      12'b101001000101 : begin
        _zz__zz_regVec_0 = regVec_2629;
      end
      12'b101001000110 : begin
        _zz__zz_regVec_0 = regVec_2630;
      end
      12'b101001000111 : begin
        _zz__zz_regVec_0 = regVec_2631;
      end
      12'b101001001000 : begin
        _zz__zz_regVec_0 = regVec_2632;
      end
      12'b101001001001 : begin
        _zz__zz_regVec_0 = regVec_2633;
      end
      12'b101001001010 : begin
        _zz__zz_regVec_0 = regVec_2634;
      end
      12'b101001001011 : begin
        _zz__zz_regVec_0 = regVec_2635;
      end
      12'b101001001100 : begin
        _zz__zz_regVec_0 = regVec_2636;
      end
      12'b101001001101 : begin
        _zz__zz_regVec_0 = regVec_2637;
      end
      12'b101001001110 : begin
        _zz__zz_regVec_0 = regVec_2638;
      end
      12'b101001001111 : begin
        _zz__zz_regVec_0 = regVec_2639;
      end
      12'b101001010000 : begin
        _zz__zz_regVec_0 = regVec_2640;
      end
      12'b101001010001 : begin
        _zz__zz_regVec_0 = regVec_2641;
      end
      12'b101001010010 : begin
        _zz__zz_regVec_0 = regVec_2642;
      end
      12'b101001010011 : begin
        _zz__zz_regVec_0 = regVec_2643;
      end
      12'b101001010100 : begin
        _zz__zz_regVec_0 = regVec_2644;
      end
      12'b101001010101 : begin
        _zz__zz_regVec_0 = regVec_2645;
      end
      12'b101001010110 : begin
        _zz__zz_regVec_0 = regVec_2646;
      end
      12'b101001010111 : begin
        _zz__zz_regVec_0 = regVec_2647;
      end
      12'b101001011000 : begin
        _zz__zz_regVec_0 = regVec_2648;
      end
      12'b101001011001 : begin
        _zz__zz_regVec_0 = regVec_2649;
      end
      12'b101001011010 : begin
        _zz__zz_regVec_0 = regVec_2650;
      end
      12'b101001011011 : begin
        _zz__zz_regVec_0 = regVec_2651;
      end
      12'b101001011100 : begin
        _zz__zz_regVec_0 = regVec_2652;
      end
      12'b101001011101 : begin
        _zz__zz_regVec_0 = regVec_2653;
      end
      12'b101001011110 : begin
        _zz__zz_regVec_0 = regVec_2654;
      end
      12'b101001011111 : begin
        _zz__zz_regVec_0 = regVec_2655;
      end
      12'b101001100000 : begin
        _zz__zz_regVec_0 = regVec_2656;
      end
      12'b101001100001 : begin
        _zz__zz_regVec_0 = regVec_2657;
      end
      12'b101001100010 : begin
        _zz__zz_regVec_0 = regVec_2658;
      end
      12'b101001100011 : begin
        _zz__zz_regVec_0 = regVec_2659;
      end
      12'b101001100100 : begin
        _zz__zz_regVec_0 = regVec_2660;
      end
      12'b101001100101 : begin
        _zz__zz_regVec_0 = regVec_2661;
      end
      12'b101001100110 : begin
        _zz__zz_regVec_0 = regVec_2662;
      end
      12'b101001100111 : begin
        _zz__zz_regVec_0 = regVec_2663;
      end
      12'b101001101000 : begin
        _zz__zz_regVec_0 = regVec_2664;
      end
      12'b101001101001 : begin
        _zz__zz_regVec_0 = regVec_2665;
      end
      12'b101001101010 : begin
        _zz__zz_regVec_0 = regVec_2666;
      end
      12'b101001101011 : begin
        _zz__zz_regVec_0 = regVec_2667;
      end
      12'b101001101100 : begin
        _zz__zz_regVec_0 = regVec_2668;
      end
      12'b101001101101 : begin
        _zz__zz_regVec_0 = regVec_2669;
      end
      12'b101001101110 : begin
        _zz__zz_regVec_0 = regVec_2670;
      end
      12'b101001101111 : begin
        _zz__zz_regVec_0 = regVec_2671;
      end
      12'b101001110000 : begin
        _zz__zz_regVec_0 = regVec_2672;
      end
      12'b101001110001 : begin
        _zz__zz_regVec_0 = regVec_2673;
      end
      12'b101001110010 : begin
        _zz__zz_regVec_0 = regVec_2674;
      end
      12'b101001110011 : begin
        _zz__zz_regVec_0 = regVec_2675;
      end
      12'b101001110100 : begin
        _zz__zz_regVec_0 = regVec_2676;
      end
      12'b101001110101 : begin
        _zz__zz_regVec_0 = regVec_2677;
      end
      12'b101001110110 : begin
        _zz__zz_regVec_0 = regVec_2678;
      end
      12'b101001110111 : begin
        _zz__zz_regVec_0 = regVec_2679;
      end
      12'b101001111000 : begin
        _zz__zz_regVec_0 = regVec_2680;
      end
      12'b101001111001 : begin
        _zz__zz_regVec_0 = regVec_2681;
      end
      12'b101001111010 : begin
        _zz__zz_regVec_0 = regVec_2682;
      end
      12'b101001111011 : begin
        _zz__zz_regVec_0 = regVec_2683;
      end
      12'b101001111100 : begin
        _zz__zz_regVec_0 = regVec_2684;
      end
      12'b101001111101 : begin
        _zz__zz_regVec_0 = regVec_2685;
      end
      12'b101001111110 : begin
        _zz__zz_regVec_0 = regVec_2686;
      end
      12'b101001111111 : begin
        _zz__zz_regVec_0 = regVec_2687;
      end
      12'b101010000000 : begin
        _zz__zz_regVec_0 = regVec_2688;
      end
      12'b101010000001 : begin
        _zz__zz_regVec_0 = regVec_2689;
      end
      12'b101010000010 : begin
        _zz__zz_regVec_0 = regVec_2690;
      end
      12'b101010000011 : begin
        _zz__zz_regVec_0 = regVec_2691;
      end
      12'b101010000100 : begin
        _zz__zz_regVec_0 = regVec_2692;
      end
      12'b101010000101 : begin
        _zz__zz_regVec_0 = regVec_2693;
      end
      12'b101010000110 : begin
        _zz__zz_regVec_0 = regVec_2694;
      end
      12'b101010000111 : begin
        _zz__zz_regVec_0 = regVec_2695;
      end
      12'b101010001000 : begin
        _zz__zz_regVec_0 = regVec_2696;
      end
      12'b101010001001 : begin
        _zz__zz_regVec_0 = regVec_2697;
      end
      12'b101010001010 : begin
        _zz__zz_regVec_0 = regVec_2698;
      end
      12'b101010001011 : begin
        _zz__zz_regVec_0 = regVec_2699;
      end
      12'b101010001100 : begin
        _zz__zz_regVec_0 = regVec_2700;
      end
      12'b101010001101 : begin
        _zz__zz_regVec_0 = regVec_2701;
      end
      12'b101010001110 : begin
        _zz__zz_regVec_0 = regVec_2702;
      end
      12'b101010001111 : begin
        _zz__zz_regVec_0 = regVec_2703;
      end
      12'b101010010000 : begin
        _zz__zz_regVec_0 = regVec_2704;
      end
      12'b101010010001 : begin
        _zz__zz_regVec_0 = regVec_2705;
      end
      12'b101010010010 : begin
        _zz__zz_regVec_0 = regVec_2706;
      end
      12'b101010010011 : begin
        _zz__zz_regVec_0 = regVec_2707;
      end
      12'b101010010100 : begin
        _zz__zz_regVec_0 = regVec_2708;
      end
      12'b101010010101 : begin
        _zz__zz_regVec_0 = regVec_2709;
      end
      12'b101010010110 : begin
        _zz__zz_regVec_0 = regVec_2710;
      end
      12'b101010010111 : begin
        _zz__zz_regVec_0 = regVec_2711;
      end
      12'b101010011000 : begin
        _zz__zz_regVec_0 = regVec_2712;
      end
      12'b101010011001 : begin
        _zz__zz_regVec_0 = regVec_2713;
      end
      12'b101010011010 : begin
        _zz__zz_regVec_0 = regVec_2714;
      end
      12'b101010011011 : begin
        _zz__zz_regVec_0 = regVec_2715;
      end
      12'b101010011100 : begin
        _zz__zz_regVec_0 = regVec_2716;
      end
      12'b101010011101 : begin
        _zz__zz_regVec_0 = regVec_2717;
      end
      12'b101010011110 : begin
        _zz__zz_regVec_0 = regVec_2718;
      end
      12'b101010011111 : begin
        _zz__zz_regVec_0 = regVec_2719;
      end
      12'b101010100000 : begin
        _zz__zz_regVec_0 = regVec_2720;
      end
      12'b101010100001 : begin
        _zz__zz_regVec_0 = regVec_2721;
      end
      12'b101010100010 : begin
        _zz__zz_regVec_0 = regVec_2722;
      end
      12'b101010100011 : begin
        _zz__zz_regVec_0 = regVec_2723;
      end
      12'b101010100100 : begin
        _zz__zz_regVec_0 = regVec_2724;
      end
      12'b101010100101 : begin
        _zz__zz_regVec_0 = regVec_2725;
      end
      12'b101010100110 : begin
        _zz__zz_regVec_0 = regVec_2726;
      end
      12'b101010100111 : begin
        _zz__zz_regVec_0 = regVec_2727;
      end
      12'b101010101000 : begin
        _zz__zz_regVec_0 = regVec_2728;
      end
      12'b101010101001 : begin
        _zz__zz_regVec_0 = regVec_2729;
      end
      12'b101010101010 : begin
        _zz__zz_regVec_0 = regVec_2730;
      end
      12'b101010101011 : begin
        _zz__zz_regVec_0 = regVec_2731;
      end
      12'b101010101100 : begin
        _zz__zz_regVec_0 = regVec_2732;
      end
      12'b101010101101 : begin
        _zz__zz_regVec_0 = regVec_2733;
      end
      12'b101010101110 : begin
        _zz__zz_regVec_0 = regVec_2734;
      end
      12'b101010101111 : begin
        _zz__zz_regVec_0 = regVec_2735;
      end
      12'b101010110000 : begin
        _zz__zz_regVec_0 = regVec_2736;
      end
      12'b101010110001 : begin
        _zz__zz_regVec_0 = regVec_2737;
      end
      12'b101010110010 : begin
        _zz__zz_regVec_0 = regVec_2738;
      end
      12'b101010110011 : begin
        _zz__zz_regVec_0 = regVec_2739;
      end
      12'b101010110100 : begin
        _zz__zz_regVec_0 = regVec_2740;
      end
      12'b101010110101 : begin
        _zz__zz_regVec_0 = regVec_2741;
      end
      12'b101010110110 : begin
        _zz__zz_regVec_0 = regVec_2742;
      end
      12'b101010110111 : begin
        _zz__zz_regVec_0 = regVec_2743;
      end
      12'b101010111000 : begin
        _zz__zz_regVec_0 = regVec_2744;
      end
      12'b101010111001 : begin
        _zz__zz_regVec_0 = regVec_2745;
      end
      12'b101010111010 : begin
        _zz__zz_regVec_0 = regVec_2746;
      end
      12'b101010111011 : begin
        _zz__zz_regVec_0 = regVec_2747;
      end
      12'b101010111100 : begin
        _zz__zz_regVec_0 = regVec_2748;
      end
      12'b101010111101 : begin
        _zz__zz_regVec_0 = regVec_2749;
      end
      12'b101010111110 : begin
        _zz__zz_regVec_0 = regVec_2750;
      end
      12'b101010111111 : begin
        _zz__zz_regVec_0 = regVec_2751;
      end
      12'b101011000000 : begin
        _zz__zz_regVec_0 = regVec_2752;
      end
      12'b101011000001 : begin
        _zz__zz_regVec_0 = regVec_2753;
      end
      12'b101011000010 : begin
        _zz__zz_regVec_0 = regVec_2754;
      end
      12'b101011000011 : begin
        _zz__zz_regVec_0 = regVec_2755;
      end
      12'b101011000100 : begin
        _zz__zz_regVec_0 = regVec_2756;
      end
      12'b101011000101 : begin
        _zz__zz_regVec_0 = regVec_2757;
      end
      12'b101011000110 : begin
        _zz__zz_regVec_0 = regVec_2758;
      end
      12'b101011000111 : begin
        _zz__zz_regVec_0 = regVec_2759;
      end
      12'b101011001000 : begin
        _zz__zz_regVec_0 = regVec_2760;
      end
      12'b101011001001 : begin
        _zz__zz_regVec_0 = regVec_2761;
      end
      12'b101011001010 : begin
        _zz__zz_regVec_0 = regVec_2762;
      end
      12'b101011001011 : begin
        _zz__zz_regVec_0 = regVec_2763;
      end
      12'b101011001100 : begin
        _zz__zz_regVec_0 = regVec_2764;
      end
      12'b101011001101 : begin
        _zz__zz_regVec_0 = regVec_2765;
      end
      12'b101011001110 : begin
        _zz__zz_regVec_0 = regVec_2766;
      end
      12'b101011001111 : begin
        _zz__zz_regVec_0 = regVec_2767;
      end
      12'b101011010000 : begin
        _zz__zz_regVec_0 = regVec_2768;
      end
      12'b101011010001 : begin
        _zz__zz_regVec_0 = regVec_2769;
      end
      12'b101011010010 : begin
        _zz__zz_regVec_0 = regVec_2770;
      end
      12'b101011010011 : begin
        _zz__zz_regVec_0 = regVec_2771;
      end
      12'b101011010100 : begin
        _zz__zz_regVec_0 = regVec_2772;
      end
      12'b101011010101 : begin
        _zz__zz_regVec_0 = regVec_2773;
      end
      12'b101011010110 : begin
        _zz__zz_regVec_0 = regVec_2774;
      end
      12'b101011010111 : begin
        _zz__zz_regVec_0 = regVec_2775;
      end
      12'b101011011000 : begin
        _zz__zz_regVec_0 = regVec_2776;
      end
      12'b101011011001 : begin
        _zz__zz_regVec_0 = regVec_2777;
      end
      12'b101011011010 : begin
        _zz__zz_regVec_0 = regVec_2778;
      end
      12'b101011011011 : begin
        _zz__zz_regVec_0 = regVec_2779;
      end
      12'b101011011100 : begin
        _zz__zz_regVec_0 = regVec_2780;
      end
      12'b101011011101 : begin
        _zz__zz_regVec_0 = regVec_2781;
      end
      12'b101011011110 : begin
        _zz__zz_regVec_0 = regVec_2782;
      end
      12'b101011011111 : begin
        _zz__zz_regVec_0 = regVec_2783;
      end
      12'b101011100000 : begin
        _zz__zz_regVec_0 = regVec_2784;
      end
      12'b101011100001 : begin
        _zz__zz_regVec_0 = regVec_2785;
      end
      12'b101011100010 : begin
        _zz__zz_regVec_0 = regVec_2786;
      end
      12'b101011100011 : begin
        _zz__zz_regVec_0 = regVec_2787;
      end
      12'b101011100100 : begin
        _zz__zz_regVec_0 = regVec_2788;
      end
      12'b101011100101 : begin
        _zz__zz_regVec_0 = regVec_2789;
      end
      12'b101011100110 : begin
        _zz__zz_regVec_0 = regVec_2790;
      end
      12'b101011100111 : begin
        _zz__zz_regVec_0 = regVec_2791;
      end
      12'b101011101000 : begin
        _zz__zz_regVec_0 = regVec_2792;
      end
      12'b101011101001 : begin
        _zz__zz_regVec_0 = regVec_2793;
      end
      12'b101011101010 : begin
        _zz__zz_regVec_0 = regVec_2794;
      end
      12'b101011101011 : begin
        _zz__zz_regVec_0 = regVec_2795;
      end
      12'b101011101100 : begin
        _zz__zz_regVec_0 = regVec_2796;
      end
      12'b101011101101 : begin
        _zz__zz_regVec_0 = regVec_2797;
      end
      12'b101011101110 : begin
        _zz__zz_regVec_0 = regVec_2798;
      end
      12'b101011101111 : begin
        _zz__zz_regVec_0 = regVec_2799;
      end
      12'b101011110000 : begin
        _zz__zz_regVec_0 = regVec_2800;
      end
      12'b101011110001 : begin
        _zz__zz_regVec_0 = regVec_2801;
      end
      12'b101011110010 : begin
        _zz__zz_regVec_0 = regVec_2802;
      end
      12'b101011110011 : begin
        _zz__zz_regVec_0 = regVec_2803;
      end
      12'b101011110100 : begin
        _zz__zz_regVec_0 = regVec_2804;
      end
      12'b101011110101 : begin
        _zz__zz_regVec_0 = regVec_2805;
      end
      12'b101011110110 : begin
        _zz__zz_regVec_0 = regVec_2806;
      end
      12'b101011110111 : begin
        _zz__zz_regVec_0 = regVec_2807;
      end
      12'b101011111000 : begin
        _zz__zz_regVec_0 = regVec_2808;
      end
      12'b101011111001 : begin
        _zz__zz_regVec_0 = regVec_2809;
      end
      12'b101011111010 : begin
        _zz__zz_regVec_0 = regVec_2810;
      end
      12'b101011111011 : begin
        _zz__zz_regVec_0 = regVec_2811;
      end
      12'b101011111100 : begin
        _zz__zz_regVec_0 = regVec_2812;
      end
      12'b101011111101 : begin
        _zz__zz_regVec_0 = regVec_2813;
      end
      12'b101011111110 : begin
        _zz__zz_regVec_0 = regVec_2814;
      end
      12'b101011111111 : begin
        _zz__zz_regVec_0 = regVec_2815;
      end
      12'b101100000000 : begin
        _zz__zz_regVec_0 = regVec_2816;
      end
      12'b101100000001 : begin
        _zz__zz_regVec_0 = regVec_2817;
      end
      12'b101100000010 : begin
        _zz__zz_regVec_0 = regVec_2818;
      end
      12'b101100000011 : begin
        _zz__zz_regVec_0 = regVec_2819;
      end
      12'b101100000100 : begin
        _zz__zz_regVec_0 = regVec_2820;
      end
      12'b101100000101 : begin
        _zz__zz_regVec_0 = regVec_2821;
      end
      12'b101100000110 : begin
        _zz__zz_regVec_0 = regVec_2822;
      end
      12'b101100000111 : begin
        _zz__zz_regVec_0 = regVec_2823;
      end
      12'b101100001000 : begin
        _zz__zz_regVec_0 = regVec_2824;
      end
      12'b101100001001 : begin
        _zz__zz_regVec_0 = regVec_2825;
      end
      12'b101100001010 : begin
        _zz__zz_regVec_0 = regVec_2826;
      end
      12'b101100001011 : begin
        _zz__zz_regVec_0 = regVec_2827;
      end
      12'b101100001100 : begin
        _zz__zz_regVec_0 = regVec_2828;
      end
      12'b101100001101 : begin
        _zz__zz_regVec_0 = regVec_2829;
      end
      12'b101100001110 : begin
        _zz__zz_regVec_0 = regVec_2830;
      end
      12'b101100001111 : begin
        _zz__zz_regVec_0 = regVec_2831;
      end
      12'b101100010000 : begin
        _zz__zz_regVec_0 = regVec_2832;
      end
      12'b101100010001 : begin
        _zz__zz_regVec_0 = regVec_2833;
      end
      12'b101100010010 : begin
        _zz__zz_regVec_0 = regVec_2834;
      end
      12'b101100010011 : begin
        _zz__zz_regVec_0 = regVec_2835;
      end
      12'b101100010100 : begin
        _zz__zz_regVec_0 = regVec_2836;
      end
      12'b101100010101 : begin
        _zz__zz_regVec_0 = regVec_2837;
      end
      12'b101100010110 : begin
        _zz__zz_regVec_0 = regVec_2838;
      end
      12'b101100010111 : begin
        _zz__zz_regVec_0 = regVec_2839;
      end
      12'b101100011000 : begin
        _zz__zz_regVec_0 = regVec_2840;
      end
      12'b101100011001 : begin
        _zz__zz_regVec_0 = regVec_2841;
      end
      12'b101100011010 : begin
        _zz__zz_regVec_0 = regVec_2842;
      end
      12'b101100011011 : begin
        _zz__zz_regVec_0 = regVec_2843;
      end
      12'b101100011100 : begin
        _zz__zz_regVec_0 = regVec_2844;
      end
      12'b101100011101 : begin
        _zz__zz_regVec_0 = regVec_2845;
      end
      12'b101100011110 : begin
        _zz__zz_regVec_0 = regVec_2846;
      end
      12'b101100011111 : begin
        _zz__zz_regVec_0 = regVec_2847;
      end
      12'b101100100000 : begin
        _zz__zz_regVec_0 = regVec_2848;
      end
      12'b101100100001 : begin
        _zz__zz_regVec_0 = regVec_2849;
      end
      12'b101100100010 : begin
        _zz__zz_regVec_0 = regVec_2850;
      end
      12'b101100100011 : begin
        _zz__zz_regVec_0 = regVec_2851;
      end
      12'b101100100100 : begin
        _zz__zz_regVec_0 = regVec_2852;
      end
      12'b101100100101 : begin
        _zz__zz_regVec_0 = regVec_2853;
      end
      12'b101100100110 : begin
        _zz__zz_regVec_0 = regVec_2854;
      end
      12'b101100100111 : begin
        _zz__zz_regVec_0 = regVec_2855;
      end
      12'b101100101000 : begin
        _zz__zz_regVec_0 = regVec_2856;
      end
      12'b101100101001 : begin
        _zz__zz_regVec_0 = regVec_2857;
      end
      12'b101100101010 : begin
        _zz__zz_regVec_0 = regVec_2858;
      end
      12'b101100101011 : begin
        _zz__zz_regVec_0 = regVec_2859;
      end
      12'b101100101100 : begin
        _zz__zz_regVec_0 = regVec_2860;
      end
      12'b101100101101 : begin
        _zz__zz_regVec_0 = regVec_2861;
      end
      12'b101100101110 : begin
        _zz__zz_regVec_0 = regVec_2862;
      end
      12'b101100101111 : begin
        _zz__zz_regVec_0 = regVec_2863;
      end
      12'b101100110000 : begin
        _zz__zz_regVec_0 = regVec_2864;
      end
      12'b101100110001 : begin
        _zz__zz_regVec_0 = regVec_2865;
      end
      12'b101100110010 : begin
        _zz__zz_regVec_0 = regVec_2866;
      end
      12'b101100110011 : begin
        _zz__zz_regVec_0 = regVec_2867;
      end
      12'b101100110100 : begin
        _zz__zz_regVec_0 = regVec_2868;
      end
      12'b101100110101 : begin
        _zz__zz_regVec_0 = regVec_2869;
      end
      12'b101100110110 : begin
        _zz__zz_regVec_0 = regVec_2870;
      end
      12'b101100110111 : begin
        _zz__zz_regVec_0 = regVec_2871;
      end
      12'b101100111000 : begin
        _zz__zz_regVec_0 = regVec_2872;
      end
      12'b101100111001 : begin
        _zz__zz_regVec_0 = regVec_2873;
      end
      12'b101100111010 : begin
        _zz__zz_regVec_0 = regVec_2874;
      end
      12'b101100111011 : begin
        _zz__zz_regVec_0 = regVec_2875;
      end
      12'b101100111100 : begin
        _zz__zz_regVec_0 = regVec_2876;
      end
      12'b101100111101 : begin
        _zz__zz_regVec_0 = regVec_2877;
      end
      12'b101100111110 : begin
        _zz__zz_regVec_0 = regVec_2878;
      end
      12'b101100111111 : begin
        _zz__zz_regVec_0 = regVec_2879;
      end
      12'b101101000000 : begin
        _zz__zz_regVec_0 = regVec_2880;
      end
      12'b101101000001 : begin
        _zz__zz_regVec_0 = regVec_2881;
      end
      12'b101101000010 : begin
        _zz__zz_regVec_0 = regVec_2882;
      end
      12'b101101000011 : begin
        _zz__zz_regVec_0 = regVec_2883;
      end
      12'b101101000100 : begin
        _zz__zz_regVec_0 = regVec_2884;
      end
      12'b101101000101 : begin
        _zz__zz_regVec_0 = regVec_2885;
      end
      12'b101101000110 : begin
        _zz__zz_regVec_0 = regVec_2886;
      end
      12'b101101000111 : begin
        _zz__zz_regVec_0 = regVec_2887;
      end
      12'b101101001000 : begin
        _zz__zz_regVec_0 = regVec_2888;
      end
      12'b101101001001 : begin
        _zz__zz_regVec_0 = regVec_2889;
      end
      12'b101101001010 : begin
        _zz__zz_regVec_0 = regVec_2890;
      end
      12'b101101001011 : begin
        _zz__zz_regVec_0 = regVec_2891;
      end
      12'b101101001100 : begin
        _zz__zz_regVec_0 = regVec_2892;
      end
      12'b101101001101 : begin
        _zz__zz_regVec_0 = regVec_2893;
      end
      12'b101101001110 : begin
        _zz__zz_regVec_0 = regVec_2894;
      end
      12'b101101001111 : begin
        _zz__zz_regVec_0 = regVec_2895;
      end
      12'b101101010000 : begin
        _zz__zz_regVec_0 = regVec_2896;
      end
      12'b101101010001 : begin
        _zz__zz_regVec_0 = regVec_2897;
      end
      12'b101101010010 : begin
        _zz__zz_regVec_0 = regVec_2898;
      end
      12'b101101010011 : begin
        _zz__zz_regVec_0 = regVec_2899;
      end
      12'b101101010100 : begin
        _zz__zz_regVec_0 = regVec_2900;
      end
      12'b101101010101 : begin
        _zz__zz_regVec_0 = regVec_2901;
      end
      12'b101101010110 : begin
        _zz__zz_regVec_0 = regVec_2902;
      end
      12'b101101010111 : begin
        _zz__zz_regVec_0 = regVec_2903;
      end
      12'b101101011000 : begin
        _zz__zz_regVec_0 = regVec_2904;
      end
      12'b101101011001 : begin
        _zz__zz_regVec_0 = regVec_2905;
      end
      12'b101101011010 : begin
        _zz__zz_regVec_0 = regVec_2906;
      end
      12'b101101011011 : begin
        _zz__zz_regVec_0 = regVec_2907;
      end
      12'b101101011100 : begin
        _zz__zz_regVec_0 = regVec_2908;
      end
      12'b101101011101 : begin
        _zz__zz_regVec_0 = regVec_2909;
      end
      12'b101101011110 : begin
        _zz__zz_regVec_0 = regVec_2910;
      end
      12'b101101011111 : begin
        _zz__zz_regVec_0 = regVec_2911;
      end
      12'b101101100000 : begin
        _zz__zz_regVec_0 = regVec_2912;
      end
      12'b101101100001 : begin
        _zz__zz_regVec_0 = regVec_2913;
      end
      12'b101101100010 : begin
        _zz__zz_regVec_0 = regVec_2914;
      end
      12'b101101100011 : begin
        _zz__zz_regVec_0 = regVec_2915;
      end
      12'b101101100100 : begin
        _zz__zz_regVec_0 = regVec_2916;
      end
      12'b101101100101 : begin
        _zz__zz_regVec_0 = regVec_2917;
      end
      12'b101101100110 : begin
        _zz__zz_regVec_0 = regVec_2918;
      end
      12'b101101100111 : begin
        _zz__zz_regVec_0 = regVec_2919;
      end
      12'b101101101000 : begin
        _zz__zz_regVec_0 = regVec_2920;
      end
      12'b101101101001 : begin
        _zz__zz_regVec_0 = regVec_2921;
      end
      12'b101101101010 : begin
        _zz__zz_regVec_0 = regVec_2922;
      end
      12'b101101101011 : begin
        _zz__zz_regVec_0 = regVec_2923;
      end
      12'b101101101100 : begin
        _zz__zz_regVec_0 = regVec_2924;
      end
      12'b101101101101 : begin
        _zz__zz_regVec_0 = regVec_2925;
      end
      12'b101101101110 : begin
        _zz__zz_regVec_0 = regVec_2926;
      end
      12'b101101101111 : begin
        _zz__zz_regVec_0 = regVec_2927;
      end
      12'b101101110000 : begin
        _zz__zz_regVec_0 = regVec_2928;
      end
      12'b101101110001 : begin
        _zz__zz_regVec_0 = regVec_2929;
      end
      12'b101101110010 : begin
        _zz__zz_regVec_0 = regVec_2930;
      end
      12'b101101110011 : begin
        _zz__zz_regVec_0 = regVec_2931;
      end
      12'b101101110100 : begin
        _zz__zz_regVec_0 = regVec_2932;
      end
      12'b101101110101 : begin
        _zz__zz_regVec_0 = regVec_2933;
      end
      12'b101101110110 : begin
        _zz__zz_regVec_0 = regVec_2934;
      end
      12'b101101110111 : begin
        _zz__zz_regVec_0 = regVec_2935;
      end
      12'b101101111000 : begin
        _zz__zz_regVec_0 = regVec_2936;
      end
      12'b101101111001 : begin
        _zz__zz_regVec_0 = regVec_2937;
      end
      12'b101101111010 : begin
        _zz__zz_regVec_0 = regVec_2938;
      end
      12'b101101111011 : begin
        _zz__zz_regVec_0 = regVec_2939;
      end
      12'b101101111100 : begin
        _zz__zz_regVec_0 = regVec_2940;
      end
      12'b101101111101 : begin
        _zz__zz_regVec_0 = regVec_2941;
      end
      12'b101101111110 : begin
        _zz__zz_regVec_0 = regVec_2942;
      end
      12'b101101111111 : begin
        _zz__zz_regVec_0 = regVec_2943;
      end
      12'b101110000000 : begin
        _zz__zz_regVec_0 = regVec_2944;
      end
      12'b101110000001 : begin
        _zz__zz_regVec_0 = regVec_2945;
      end
      12'b101110000010 : begin
        _zz__zz_regVec_0 = regVec_2946;
      end
      12'b101110000011 : begin
        _zz__zz_regVec_0 = regVec_2947;
      end
      12'b101110000100 : begin
        _zz__zz_regVec_0 = regVec_2948;
      end
      12'b101110000101 : begin
        _zz__zz_regVec_0 = regVec_2949;
      end
      12'b101110000110 : begin
        _zz__zz_regVec_0 = regVec_2950;
      end
      12'b101110000111 : begin
        _zz__zz_regVec_0 = regVec_2951;
      end
      12'b101110001000 : begin
        _zz__zz_regVec_0 = regVec_2952;
      end
      12'b101110001001 : begin
        _zz__zz_regVec_0 = regVec_2953;
      end
      12'b101110001010 : begin
        _zz__zz_regVec_0 = regVec_2954;
      end
      12'b101110001011 : begin
        _zz__zz_regVec_0 = regVec_2955;
      end
      12'b101110001100 : begin
        _zz__zz_regVec_0 = regVec_2956;
      end
      12'b101110001101 : begin
        _zz__zz_regVec_0 = regVec_2957;
      end
      12'b101110001110 : begin
        _zz__zz_regVec_0 = regVec_2958;
      end
      12'b101110001111 : begin
        _zz__zz_regVec_0 = regVec_2959;
      end
      12'b101110010000 : begin
        _zz__zz_regVec_0 = regVec_2960;
      end
      12'b101110010001 : begin
        _zz__zz_regVec_0 = regVec_2961;
      end
      12'b101110010010 : begin
        _zz__zz_regVec_0 = regVec_2962;
      end
      12'b101110010011 : begin
        _zz__zz_regVec_0 = regVec_2963;
      end
      12'b101110010100 : begin
        _zz__zz_regVec_0 = regVec_2964;
      end
      12'b101110010101 : begin
        _zz__zz_regVec_0 = regVec_2965;
      end
      12'b101110010110 : begin
        _zz__zz_regVec_0 = regVec_2966;
      end
      12'b101110010111 : begin
        _zz__zz_regVec_0 = regVec_2967;
      end
      12'b101110011000 : begin
        _zz__zz_regVec_0 = regVec_2968;
      end
      12'b101110011001 : begin
        _zz__zz_regVec_0 = regVec_2969;
      end
      12'b101110011010 : begin
        _zz__zz_regVec_0 = regVec_2970;
      end
      12'b101110011011 : begin
        _zz__zz_regVec_0 = regVec_2971;
      end
      12'b101110011100 : begin
        _zz__zz_regVec_0 = regVec_2972;
      end
      12'b101110011101 : begin
        _zz__zz_regVec_0 = regVec_2973;
      end
      12'b101110011110 : begin
        _zz__zz_regVec_0 = regVec_2974;
      end
      12'b101110011111 : begin
        _zz__zz_regVec_0 = regVec_2975;
      end
      12'b101110100000 : begin
        _zz__zz_regVec_0 = regVec_2976;
      end
      12'b101110100001 : begin
        _zz__zz_regVec_0 = regVec_2977;
      end
      12'b101110100010 : begin
        _zz__zz_regVec_0 = regVec_2978;
      end
      12'b101110100011 : begin
        _zz__zz_regVec_0 = regVec_2979;
      end
      12'b101110100100 : begin
        _zz__zz_regVec_0 = regVec_2980;
      end
      12'b101110100101 : begin
        _zz__zz_regVec_0 = regVec_2981;
      end
      12'b101110100110 : begin
        _zz__zz_regVec_0 = regVec_2982;
      end
      12'b101110100111 : begin
        _zz__zz_regVec_0 = regVec_2983;
      end
      12'b101110101000 : begin
        _zz__zz_regVec_0 = regVec_2984;
      end
      12'b101110101001 : begin
        _zz__zz_regVec_0 = regVec_2985;
      end
      12'b101110101010 : begin
        _zz__zz_regVec_0 = regVec_2986;
      end
      12'b101110101011 : begin
        _zz__zz_regVec_0 = regVec_2987;
      end
      12'b101110101100 : begin
        _zz__zz_regVec_0 = regVec_2988;
      end
      12'b101110101101 : begin
        _zz__zz_regVec_0 = regVec_2989;
      end
      12'b101110101110 : begin
        _zz__zz_regVec_0 = regVec_2990;
      end
      12'b101110101111 : begin
        _zz__zz_regVec_0 = regVec_2991;
      end
      12'b101110110000 : begin
        _zz__zz_regVec_0 = regVec_2992;
      end
      12'b101110110001 : begin
        _zz__zz_regVec_0 = regVec_2993;
      end
      12'b101110110010 : begin
        _zz__zz_regVec_0 = regVec_2994;
      end
      12'b101110110011 : begin
        _zz__zz_regVec_0 = regVec_2995;
      end
      12'b101110110100 : begin
        _zz__zz_regVec_0 = regVec_2996;
      end
      12'b101110110101 : begin
        _zz__zz_regVec_0 = regVec_2997;
      end
      12'b101110110110 : begin
        _zz__zz_regVec_0 = regVec_2998;
      end
      12'b101110110111 : begin
        _zz__zz_regVec_0 = regVec_2999;
      end
      12'b101110111000 : begin
        _zz__zz_regVec_0 = regVec_3000;
      end
      12'b101110111001 : begin
        _zz__zz_regVec_0 = regVec_3001;
      end
      12'b101110111010 : begin
        _zz__zz_regVec_0 = regVec_3002;
      end
      12'b101110111011 : begin
        _zz__zz_regVec_0 = regVec_3003;
      end
      12'b101110111100 : begin
        _zz__zz_regVec_0 = regVec_3004;
      end
      12'b101110111101 : begin
        _zz__zz_regVec_0 = regVec_3005;
      end
      12'b101110111110 : begin
        _zz__zz_regVec_0 = regVec_3006;
      end
      12'b101110111111 : begin
        _zz__zz_regVec_0 = regVec_3007;
      end
      12'b101111000000 : begin
        _zz__zz_regVec_0 = regVec_3008;
      end
      12'b101111000001 : begin
        _zz__zz_regVec_0 = regVec_3009;
      end
      12'b101111000010 : begin
        _zz__zz_regVec_0 = regVec_3010;
      end
      12'b101111000011 : begin
        _zz__zz_regVec_0 = regVec_3011;
      end
      12'b101111000100 : begin
        _zz__zz_regVec_0 = regVec_3012;
      end
      12'b101111000101 : begin
        _zz__zz_regVec_0 = regVec_3013;
      end
      12'b101111000110 : begin
        _zz__zz_regVec_0 = regVec_3014;
      end
      12'b101111000111 : begin
        _zz__zz_regVec_0 = regVec_3015;
      end
      12'b101111001000 : begin
        _zz__zz_regVec_0 = regVec_3016;
      end
      12'b101111001001 : begin
        _zz__zz_regVec_0 = regVec_3017;
      end
      12'b101111001010 : begin
        _zz__zz_regVec_0 = regVec_3018;
      end
      12'b101111001011 : begin
        _zz__zz_regVec_0 = regVec_3019;
      end
      12'b101111001100 : begin
        _zz__zz_regVec_0 = regVec_3020;
      end
      12'b101111001101 : begin
        _zz__zz_regVec_0 = regVec_3021;
      end
      12'b101111001110 : begin
        _zz__zz_regVec_0 = regVec_3022;
      end
      12'b101111001111 : begin
        _zz__zz_regVec_0 = regVec_3023;
      end
      12'b101111010000 : begin
        _zz__zz_regVec_0 = regVec_3024;
      end
      12'b101111010001 : begin
        _zz__zz_regVec_0 = regVec_3025;
      end
      12'b101111010010 : begin
        _zz__zz_regVec_0 = regVec_3026;
      end
      12'b101111010011 : begin
        _zz__zz_regVec_0 = regVec_3027;
      end
      12'b101111010100 : begin
        _zz__zz_regVec_0 = regVec_3028;
      end
      12'b101111010101 : begin
        _zz__zz_regVec_0 = regVec_3029;
      end
      12'b101111010110 : begin
        _zz__zz_regVec_0 = regVec_3030;
      end
      12'b101111010111 : begin
        _zz__zz_regVec_0 = regVec_3031;
      end
      12'b101111011000 : begin
        _zz__zz_regVec_0 = regVec_3032;
      end
      12'b101111011001 : begin
        _zz__zz_regVec_0 = regVec_3033;
      end
      12'b101111011010 : begin
        _zz__zz_regVec_0 = regVec_3034;
      end
      12'b101111011011 : begin
        _zz__zz_regVec_0 = regVec_3035;
      end
      12'b101111011100 : begin
        _zz__zz_regVec_0 = regVec_3036;
      end
      12'b101111011101 : begin
        _zz__zz_regVec_0 = regVec_3037;
      end
      12'b101111011110 : begin
        _zz__zz_regVec_0 = regVec_3038;
      end
      12'b101111011111 : begin
        _zz__zz_regVec_0 = regVec_3039;
      end
      12'b101111100000 : begin
        _zz__zz_regVec_0 = regVec_3040;
      end
      12'b101111100001 : begin
        _zz__zz_regVec_0 = regVec_3041;
      end
      12'b101111100010 : begin
        _zz__zz_regVec_0 = regVec_3042;
      end
      12'b101111100011 : begin
        _zz__zz_regVec_0 = regVec_3043;
      end
      12'b101111100100 : begin
        _zz__zz_regVec_0 = regVec_3044;
      end
      12'b101111100101 : begin
        _zz__zz_regVec_0 = regVec_3045;
      end
      12'b101111100110 : begin
        _zz__zz_regVec_0 = regVec_3046;
      end
      12'b101111100111 : begin
        _zz__zz_regVec_0 = regVec_3047;
      end
      12'b101111101000 : begin
        _zz__zz_regVec_0 = regVec_3048;
      end
      12'b101111101001 : begin
        _zz__zz_regVec_0 = regVec_3049;
      end
      12'b101111101010 : begin
        _zz__zz_regVec_0 = regVec_3050;
      end
      12'b101111101011 : begin
        _zz__zz_regVec_0 = regVec_3051;
      end
      12'b101111101100 : begin
        _zz__zz_regVec_0 = regVec_3052;
      end
      12'b101111101101 : begin
        _zz__zz_regVec_0 = regVec_3053;
      end
      12'b101111101110 : begin
        _zz__zz_regVec_0 = regVec_3054;
      end
      12'b101111101111 : begin
        _zz__zz_regVec_0 = regVec_3055;
      end
      12'b101111110000 : begin
        _zz__zz_regVec_0 = regVec_3056;
      end
      12'b101111110001 : begin
        _zz__zz_regVec_0 = regVec_3057;
      end
      12'b101111110010 : begin
        _zz__zz_regVec_0 = regVec_3058;
      end
      12'b101111110011 : begin
        _zz__zz_regVec_0 = regVec_3059;
      end
      12'b101111110100 : begin
        _zz__zz_regVec_0 = regVec_3060;
      end
      12'b101111110101 : begin
        _zz__zz_regVec_0 = regVec_3061;
      end
      12'b101111110110 : begin
        _zz__zz_regVec_0 = regVec_3062;
      end
      12'b101111110111 : begin
        _zz__zz_regVec_0 = regVec_3063;
      end
      12'b101111111000 : begin
        _zz__zz_regVec_0 = regVec_3064;
      end
      12'b101111111001 : begin
        _zz__zz_regVec_0 = regVec_3065;
      end
      12'b101111111010 : begin
        _zz__zz_regVec_0 = regVec_3066;
      end
      12'b101111111011 : begin
        _zz__zz_regVec_0 = regVec_3067;
      end
      12'b101111111100 : begin
        _zz__zz_regVec_0 = regVec_3068;
      end
      12'b101111111101 : begin
        _zz__zz_regVec_0 = regVec_3069;
      end
      12'b101111111110 : begin
        _zz__zz_regVec_0 = regVec_3070;
      end
      12'b101111111111 : begin
        _zz__zz_regVec_0 = regVec_3071;
      end
      12'b110000000000 : begin
        _zz__zz_regVec_0 = regVec_3072;
      end
      12'b110000000001 : begin
        _zz__zz_regVec_0 = regVec_3073;
      end
      12'b110000000010 : begin
        _zz__zz_regVec_0 = regVec_3074;
      end
      12'b110000000011 : begin
        _zz__zz_regVec_0 = regVec_3075;
      end
      12'b110000000100 : begin
        _zz__zz_regVec_0 = regVec_3076;
      end
      12'b110000000101 : begin
        _zz__zz_regVec_0 = regVec_3077;
      end
      12'b110000000110 : begin
        _zz__zz_regVec_0 = regVec_3078;
      end
      12'b110000000111 : begin
        _zz__zz_regVec_0 = regVec_3079;
      end
      12'b110000001000 : begin
        _zz__zz_regVec_0 = regVec_3080;
      end
      12'b110000001001 : begin
        _zz__zz_regVec_0 = regVec_3081;
      end
      12'b110000001010 : begin
        _zz__zz_regVec_0 = regVec_3082;
      end
      12'b110000001011 : begin
        _zz__zz_regVec_0 = regVec_3083;
      end
      12'b110000001100 : begin
        _zz__zz_regVec_0 = regVec_3084;
      end
      12'b110000001101 : begin
        _zz__zz_regVec_0 = regVec_3085;
      end
      12'b110000001110 : begin
        _zz__zz_regVec_0 = regVec_3086;
      end
      12'b110000001111 : begin
        _zz__zz_regVec_0 = regVec_3087;
      end
      12'b110000010000 : begin
        _zz__zz_regVec_0 = regVec_3088;
      end
      12'b110000010001 : begin
        _zz__zz_regVec_0 = regVec_3089;
      end
      12'b110000010010 : begin
        _zz__zz_regVec_0 = regVec_3090;
      end
      12'b110000010011 : begin
        _zz__zz_regVec_0 = regVec_3091;
      end
      12'b110000010100 : begin
        _zz__zz_regVec_0 = regVec_3092;
      end
      12'b110000010101 : begin
        _zz__zz_regVec_0 = regVec_3093;
      end
      12'b110000010110 : begin
        _zz__zz_regVec_0 = regVec_3094;
      end
      12'b110000010111 : begin
        _zz__zz_regVec_0 = regVec_3095;
      end
      12'b110000011000 : begin
        _zz__zz_regVec_0 = regVec_3096;
      end
      12'b110000011001 : begin
        _zz__zz_regVec_0 = regVec_3097;
      end
      12'b110000011010 : begin
        _zz__zz_regVec_0 = regVec_3098;
      end
      12'b110000011011 : begin
        _zz__zz_regVec_0 = regVec_3099;
      end
      12'b110000011100 : begin
        _zz__zz_regVec_0 = regVec_3100;
      end
      12'b110000011101 : begin
        _zz__zz_regVec_0 = regVec_3101;
      end
      12'b110000011110 : begin
        _zz__zz_regVec_0 = regVec_3102;
      end
      12'b110000011111 : begin
        _zz__zz_regVec_0 = regVec_3103;
      end
      12'b110000100000 : begin
        _zz__zz_regVec_0 = regVec_3104;
      end
      12'b110000100001 : begin
        _zz__zz_regVec_0 = regVec_3105;
      end
      12'b110000100010 : begin
        _zz__zz_regVec_0 = regVec_3106;
      end
      12'b110000100011 : begin
        _zz__zz_regVec_0 = regVec_3107;
      end
      12'b110000100100 : begin
        _zz__zz_regVec_0 = regVec_3108;
      end
      12'b110000100101 : begin
        _zz__zz_regVec_0 = regVec_3109;
      end
      12'b110000100110 : begin
        _zz__zz_regVec_0 = regVec_3110;
      end
      12'b110000100111 : begin
        _zz__zz_regVec_0 = regVec_3111;
      end
      12'b110000101000 : begin
        _zz__zz_regVec_0 = regVec_3112;
      end
      12'b110000101001 : begin
        _zz__zz_regVec_0 = regVec_3113;
      end
      12'b110000101010 : begin
        _zz__zz_regVec_0 = regVec_3114;
      end
      12'b110000101011 : begin
        _zz__zz_regVec_0 = regVec_3115;
      end
      12'b110000101100 : begin
        _zz__zz_regVec_0 = regVec_3116;
      end
      12'b110000101101 : begin
        _zz__zz_regVec_0 = regVec_3117;
      end
      12'b110000101110 : begin
        _zz__zz_regVec_0 = regVec_3118;
      end
      12'b110000101111 : begin
        _zz__zz_regVec_0 = regVec_3119;
      end
      12'b110000110000 : begin
        _zz__zz_regVec_0 = regVec_3120;
      end
      12'b110000110001 : begin
        _zz__zz_regVec_0 = regVec_3121;
      end
      12'b110000110010 : begin
        _zz__zz_regVec_0 = regVec_3122;
      end
      12'b110000110011 : begin
        _zz__zz_regVec_0 = regVec_3123;
      end
      12'b110000110100 : begin
        _zz__zz_regVec_0 = regVec_3124;
      end
      12'b110000110101 : begin
        _zz__zz_regVec_0 = regVec_3125;
      end
      12'b110000110110 : begin
        _zz__zz_regVec_0 = regVec_3126;
      end
      12'b110000110111 : begin
        _zz__zz_regVec_0 = regVec_3127;
      end
      12'b110000111000 : begin
        _zz__zz_regVec_0 = regVec_3128;
      end
      12'b110000111001 : begin
        _zz__zz_regVec_0 = regVec_3129;
      end
      12'b110000111010 : begin
        _zz__zz_regVec_0 = regVec_3130;
      end
      12'b110000111011 : begin
        _zz__zz_regVec_0 = regVec_3131;
      end
      12'b110000111100 : begin
        _zz__zz_regVec_0 = regVec_3132;
      end
      12'b110000111101 : begin
        _zz__zz_regVec_0 = regVec_3133;
      end
      12'b110000111110 : begin
        _zz__zz_regVec_0 = regVec_3134;
      end
      12'b110000111111 : begin
        _zz__zz_regVec_0 = regVec_3135;
      end
      12'b110001000000 : begin
        _zz__zz_regVec_0 = regVec_3136;
      end
      12'b110001000001 : begin
        _zz__zz_regVec_0 = regVec_3137;
      end
      12'b110001000010 : begin
        _zz__zz_regVec_0 = regVec_3138;
      end
      12'b110001000011 : begin
        _zz__zz_regVec_0 = regVec_3139;
      end
      12'b110001000100 : begin
        _zz__zz_regVec_0 = regVec_3140;
      end
      12'b110001000101 : begin
        _zz__zz_regVec_0 = regVec_3141;
      end
      12'b110001000110 : begin
        _zz__zz_regVec_0 = regVec_3142;
      end
      12'b110001000111 : begin
        _zz__zz_regVec_0 = regVec_3143;
      end
      12'b110001001000 : begin
        _zz__zz_regVec_0 = regVec_3144;
      end
      12'b110001001001 : begin
        _zz__zz_regVec_0 = regVec_3145;
      end
      12'b110001001010 : begin
        _zz__zz_regVec_0 = regVec_3146;
      end
      12'b110001001011 : begin
        _zz__zz_regVec_0 = regVec_3147;
      end
      12'b110001001100 : begin
        _zz__zz_regVec_0 = regVec_3148;
      end
      12'b110001001101 : begin
        _zz__zz_regVec_0 = regVec_3149;
      end
      12'b110001001110 : begin
        _zz__zz_regVec_0 = regVec_3150;
      end
      12'b110001001111 : begin
        _zz__zz_regVec_0 = regVec_3151;
      end
      12'b110001010000 : begin
        _zz__zz_regVec_0 = regVec_3152;
      end
      12'b110001010001 : begin
        _zz__zz_regVec_0 = regVec_3153;
      end
      12'b110001010010 : begin
        _zz__zz_regVec_0 = regVec_3154;
      end
      12'b110001010011 : begin
        _zz__zz_regVec_0 = regVec_3155;
      end
      12'b110001010100 : begin
        _zz__zz_regVec_0 = regVec_3156;
      end
      12'b110001010101 : begin
        _zz__zz_regVec_0 = regVec_3157;
      end
      12'b110001010110 : begin
        _zz__zz_regVec_0 = regVec_3158;
      end
      12'b110001010111 : begin
        _zz__zz_regVec_0 = regVec_3159;
      end
      12'b110001011000 : begin
        _zz__zz_regVec_0 = regVec_3160;
      end
      12'b110001011001 : begin
        _zz__zz_regVec_0 = regVec_3161;
      end
      12'b110001011010 : begin
        _zz__zz_regVec_0 = regVec_3162;
      end
      12'b110001011011 : begin
        _zz__zz_regVec_0 = regVec_3163;
      end
      12'b110001011100 : begin
        _zz__zz_regVec_0 = regVec_3164;
      end
      12'b110001011101 : begin
        _zz__zz_regVec_0 = regVec_3165;
      end
      12'b110001011110 : begin
        _zz__zz_regVec_0 = regVec_3166;
      end
      12'b110001011111 : begin
        _zz__zz_regVec_0 = regVec_3167;
      end
      12'b110001100000 : begin
        _zz__zz_regVec_0 = regVec_3168;
      end
      12'b110001100001 : begin
        _zz__zz_regVec_0 = regVec_3169;
      end
      12'b110001100010 : begin
        _zz__zz_regVec_0 = regVec_3170;
      end
      12'b110001100011 : begin
        _zz__zz_regVec_0 = regVec_3171;
      end
      12'b110001100100 : begin
        _zz__zz_regVec_0 = regVec_3172;
      end
      12'b110001100101 : begin
        _zz__zz_regVec_0 = regVec_3173;
      end
      12'b110001100110 : begin
        _zz__zz_regVec_0 = regVec_3174;
      end
      12'b110001100111 : begin
        _zz__zz_regVec_0 = regVec_3175;
      end
      12'b110001101000 : begin
        _zz__zz_regVec_0 = regVec_3176;
      end
      12'b110001101001 : begin
        _zz__zz_regVec_0 = regVec_3177;
      end
      12'b110001101010 : begin
        _zz__zz_regVec_0 = regVec_3178;
      end
      12'b110001101011 : begin
        _zz__zz_regVec_0 = regVec_3179;
      end
      12'b110001101100 : begin
        _zz__zz_regVec_0 = regVec_3180;
      end
      12'b110001101101 : begin
        _zz__zz_regVec_0 = regVec_3181;
      end
      12'b110001101110 : begin
        _zz__zz_regVec_0 = regVec_3182;
      end
      12'b110001101111 : begin
        _zz__zz_regVec_0 = regVec_3183;
      end
      12'b110001110000 : begin
        _zz__zz_regVec_0 = regVec_3184;
      end
      12'b110001110001 : begin
        _zz__zz_regVec_0 = regVec_3185;
      end
      12'b110001110010 : begin
        _zz__zz_regVec_0 = regVec_3186;
      end
      12'b110001110011 : begin
        _zz__zz_regVec_0 = regVec_3187;
      end
      12'b110001110100 : begin
        _zz__zz_regVec_0 = regVec_3188;
      end
      12'b110001110101 : begin
        _zz__zz_regVec_0 = regVec_3189;
      end
      12'b110001110110 : begin
        _zz__zz_regVec_0 = regVec_3190;
      end
      12'b110001110111 : begin
        _zz__zz_regVec_0 = regVec_3191;
      end
      12'b110001111000 : begin
        _zz__zz_regVec_0 = regVec_3192;
      end
      12'b110001111001 : begin
        _zz__zz_regVec_0 = regVec_3193;
      end
      12'b110001111010 : begin
        _zz__zz_regVec_0 = regVec_3194;
      end
      12'b110001111011 : begin
        _zz__zz_regVec_0 = regVec_3195;
      end
      12'b110001111100 : begin
        _zz__zz_regVec_0 = regVec_3196;
      end
      12'b110001111101 : begin
        _zz__zz_regVec_0 = regVec_3197;
      end
      12'b110001111110 : begin
        _zz__zz_regVec_0 = regVec_3198;
      end
      12'b110001111111 : begin
        _zz__zz_regVec_0 = regVec_3199;
      end
      12'b110010000000 : begin
        _zz__zz_regVec_0 = regVec_3200;
      end
      12'b110010000001 : begin
        _zz__zz_regVec_0 = regVec_3201;
      end
      12'b110010000010 : begin
        _zz__zz_regVec_0 = regVec_3202;
      end
      12'b110010000011 : begin
        _zz__zz_regVec_0 = regVec_3203;
      end
      12'b110010000100 : begin
        _zz__zz_regVec_0 = regVec_3204;
      end
      12'b110010000101 : begin
        _zz__zz_regVec_0 = regVec_3205;
      end
      12'b110010000110 : begin
        _zz__zz_regVec_0 = regVec_3206;
      end
      12'b110010000111 : begin
        _zz__zz_regVec_0 = regVec_3207;
      end
      12'b110010001000 : begin
        _zz__zz_regVec_0 = regVec_3208;
      end
      12'b110010001001 : begin
        _zz__zz_regVec_0 = regVec_3209;
      end
      12'b110010001010 : begin
        _zz__zz_regVec_0 = regVec_3210;
      end
      12'b110010001011 : begin
        _zz__zz_regVec_0 = regVec_3211;
      end
      12'b110010001100 : begin
        _zz__zz_regVec_0 = regVec_3212;
      end
      12'b110010001101 : begin
        _zz__zz_regVec_0 = regVec_3213;
      end
      12'b110010001110 : begin
        _zz__zz_regVec_0 = regVec_3214;
      end
      12'b110010001111 : begin
        _zz__zz_regVec_0 = regVec_3215;
      end
      12'b110010010000 : begin
        _zz__zz_regVec_0 = regVec_3216;
      end
      12'b110010010001 : begin
        _zz__zz_regVec_0 = regVec_3217;
      end
      12'b110010010010 : begin
        _zz__zz_regVec_0 = regVec_3218;
      end
      12'b110010010011 : begin
        _zz__zz_regVec_0 = regVec_3219;
      end
      12'b110010010100 : begin
        _zz__zz_regVec_0 = regVec_3220;
      end
      12'b110010010101 : begin
        _zz__zz_regVec_0 = regVec_3221;
      end
      12'b110010010110 : begin
        _zz__zz_regVec_0 = regVec_3222;
      end
      12'b110010010111 : begin
        _zz__zz_regVec_0 = regVec_3223;
      end
      12'b110010011000 : begin
        _zz__zz_regVec_0 = regVec_3224;
      end
      12'b110010011001 : begin
        _zz__zz_regVec_0 = regVec_3225;
      end
      12'b110010011010 : begin
        _zz__zz_regVec_0 = regVec_3226;
      end
      12'b110010011011 : begin
        _zz__zz_regVec_0 = regVec_3227;
      end
      12'b110010011100 : begin
        _zz__zz_regVec_0 = regVec_3228;
      end
      12'b110010011101 : begin
        _zz__zz_regVec_0 = regVec_3229;
      end
      12'b110010011110 : begin
        _zz__zz_regVec_0 = regVec_3230;
      end
      12'b110010011111 : begin
        _zz__zz_regVec_0 = regVec_3231;
      end
      12'b110010100000 : begin
        _zz__zz_regVec_0 = regVec_3232;
      end
      12'b110010100001 : begin
        _zz__zz_regVec_0 = regVec_3233;
      end
      12'b110010100010 : begin
        _zz__zz_regVec_0 = regVec_3234;
      end
      12'b110010100011 : begin
        _zz__zz_regVec_0 = regVec_3235;
      end
      12'b110010100100 : begin
        _zz__zz_regVec_0 = regVec_3236;
      end
      12'b110010100101 : begin
        _zz__zz_regVec_0 = regVec_3237;
      end
      12'b110010100110 : begin
        _zz__zz_regVec_0 = regVec_3238;
      end
      12'b110010100111 : begin
        _zz__zz_regVec_0 = regVec_3239;
      end
      12'b110010101000 : begin
        _zz__zz_regVec_0 = regVec_3240;
      end
      12'b110010101001 : begin
        _zz__zz_regVec_0 = regVec_3241;
      end
      12'b110010101010 : begin
        _zz__zz_regVec_0 = regVec_3242;
      end
      12'b110010101011 : begin
        _zz__zz_regVec_0 = regVec_3243;
      end
      12'b110010101100 : begin
        _zz__zz_regVec_0 = regVec_3244;
      end
      12'b110010101101 : begin
        _zz__zz_regVec_0 = regVec_3245;
      end
      12'b110010101110 : begin
        _zz__zz_regVec_0 = regVec_3246;
      end
      12'b110010101111 : begin
        _zz__zz_regVec_0 = regVec_3247;
      end
      12'b110010110000 : begin
        _zz__zz_regVec_0 = regVec_3248;
      end
      12'b110010110001 : begin
        _zz__zz_regVec_0 = regVec_3249;
      end
      12'b110010110010 : begin
        _zz__zz_regVec_0 = regVec_3250;
      end
      12'b110010110011 : begin
        _zz__zz_regVec_0 = regVec_3251;
      end
      12'b110010110100 : begin
        _zz__zz_regVec_0 = regVec_3252;
      end
      12'b110010110101 : begin
        _zz__zz_regVec_0 = regVec_3253;
      end
      12'b110010110110 : begin
        _zz__zz_regVec_0 = regVec_3254;
      end
      12'b110010110111 : begin
        _zz__zz_regVec_0 = regVec_3255;
      end
      12'b110010111000 : begin
        _zz__zz_regVec_0 = regVec_3256;
      end
      12'b110010111001 : begin
        _zz__zz_regVec_0 = regVec_3257;
      end
      12'b110010111010 : begin
        _zz__zz_regVec_0 = regVec_3258;
      end
      12'b110010111011 : begin
        _zz__zz_regVec_0 = regVec_3259;
      end
      12'b110010111100 : begin
        _zz__zz_regVec_0 = regVec_3260;
      end
      12'b110010111101 : begin
        _zz__zz_regVec_0 = regVec_3261;
      end
      12'b110010111110 : begin
        _zz__zz_regVec_0 = regVec_3262;
      end
      12'b110010111111 : begin
        _zz__zz_regVec_0 = regVec_3263;
      end
      12'b110011000000 : begin
        _zz__zz_regVec_0 = regVec_3264;
      end
      12'b110011000001 : begin
        _zz__zz_regVec_0 = regVec_3265;
      end
      12'b110011000010 : begin
        _zz__zz_regVec_0 = regVec_3266;
      end
      12'b110011000011 : begin
        _zz__zz_regVec_0 = regVec_3267;
      end
      12'b110011000100 : begin
        _zz__zz_regVec_0 = regVec_3268;
      end
      12'b110011000101 : begin
        _zz__zz_regVec_0 = regVec_3269;
      end
      12'b110011000110 : begin
        _zz__zz_regVec_0 = regVec_3270;
      end
      12'b110011000111 : begin
        _zz__zz_regVec_0 = regVec_3271;
      end
      12'b110011001000 : begin
        _zz__zz_regVec_0 = regVec_3272;
      end
      12'b110011001001 : begin
        _zz__zz_regVec_0 = regVec_3273;
      end
      12'b110011001010 : begin
        _zz__zz_regVec_0 = regVec_3274;
      end
      12'b110011001011 : begin
        _zz__zz_regVec_0 = regVec_3275;
      end
      12'b110011001100 : begin
        _zz__zz_regVec_0 = regVec_3276;
      end
      12'b110011001101 : begin
        _zz__zz_regVec_0 = regVec_3277;
      end
      12'b110011001110 : begin
        _zz__zz_regVec_0 = regVec_3278;
      end
      12'b110011001111 : begin
        _zz__zz_regVec_0 = regVec_3279;
      end
      12'b110011010000 : begin
        _zz__zz_regVec_0 = regVec_3280;
      end
      12'b110011010001 : begin
        _zz__zz_regVec_0 = regVec_3281;
      end
      12'b110011010010 : begin
        _zz__zz_regVec_0 = regVec_3282;
      end
      12'b110011010011 : begin
        _zz__zz_regVec_0 = regVec_3283;
      end
      12'b110011010100 : begin
        _zz__zz_regVec_0 = regVec_3284;
      end
      12'b110011010101 : begin
        _zz__zz_regVec_0 = regVec_3285;
      end
      12'b110011010110 : begin
        _zz__zz_regVec_0 = regVec_3286;
      end
      12'b110011010111 : begin
        _zz__zz_regVec_0 = regVec_3287;
      end
      12'b110011011000 : begin
        _zz__zz_regVec_0 = regVec_3288;
      end
      12'b110011011001 : begin
        _zz__zz_regVec_0 = regVec_3289;
      end
      12'b110011011010 : begin
        _zz__zz_regVec_0 = regVec_3290;
      end
      12'b110011011011 : begin
        _zz__zz_regVec_0 = regVec_3291;
      end
      12'b110011011100 : begin
        _zz__zz_regVec_0 = regVec_3292;
      end
      12'b110011011101 : begin
        _zz__zz_regVec_0 = regVec_3293;
      end
      12'b110011011110 : begin
        _zz__zz_regVec_0 = regVec_3294;
      end
      12'b110011011111 : begin
        _zz__zz_regVec_0 = regVec_3295;
      end
      12'b110011100000 : begin
        _zz__zz_regVec_0 = regVec_3296;
      end
      12'b110011100001 : begin
        _zz__zz_regVec_0 = regVec_3297;
      end
      12'b110011100010 : begin
        _zz__zz_regVec_0 = regVec_3298;
      end
      12'b110011100011 : begin
        _zz__zz_regVec_0 = regVec_3299;
      end
      12'b110011100100 : begin
        _zz__zz_regVec_0 = regVec_3300;
      end
      12'b110011100101 : begin
        _zz__zz_regVec_0 = regVec_3301;
      end
      12'b110011100110 : begin
        _zz__zz_regVec_0 = regVec_3302;
      end
      12'b110011100111 : begin
        _zz__zz_regVec_0 = regVec_3303;
      end
      12'b110011101000 : begin
        _zz__zz_regVec_0 = regVec_3304;
      end
      12'b110011101001 : begin
        _zz__zz_regVec_0 = regVec_3305;
      end
      12'b110011101010 : begin
        _zz__zz_regVec_0 = regVec_3306;
      end
      12'b110011101011 : begin
        _zz__zz_regVec_0 = regVec_3307;
      end
      12'b110011101100 : begin
        _zz__zz_regVec_0 = regVec_3308;
      end
      12'b110011101101 : begin
        _zz__zz_regVec_0 = regVec_3309;
      end
      12'b110011101110 : begin
        _zz__zz_regVec_0 = regVec_3310;
      end
      12'b110011101111 : begin
        _zz__zz_regVec_0 = regVec_3311;
      end
      12'b110011110000 : begin
        _zz__zz_regVec_0 = regVec_3312;
      end
      12'b110011110001 : begin
        _zz__zz_regVec_0 = regVec_3313;
      end
      12'b110011110010 : begin
        _zz__zz_regVec_0 = regVec_3314;
      end
      12'b110011110011 : begin
        _zz__zz_regVec_0 = regVec_3315;
      end
      12'b110011110100 : begin
        _zz__zz_regVec_0 = regVec_3316;
      end
      12'b110011110101 : begin
        _zz__zz_regVec_0 = regVec_3317;
      end
      12'b110011110110 : begin
        _zz__zz_regVec_0 = regVec_3318;
      end
      12'b110011110111 : begin
        _zz__zz_regVec_0 = regVec_3319;
      end
      12'b110011111000 : begin
        _zz__zz_regVec_0 = regVec_3320;
      end
      12'b110011111001 : begin
        _zz__zz_regVec_0 = regVec_3321;
      end
      12'b110011111010 : begin
        _zz__zz_regVec_0 = regVec_3322;
      end
      12'b110011111011 : begin
        _zz__zz_regVec_0 = regVec_3323;
      end
      12'b110011111100 : begin
        _zz__zz_regVec_0 = regVec_3324;
      end
      12'b110011111101 : begin
        _zz__zz_regVec_0 = regVec_3325;
      end
      12'b110011111110 : begin
        _zz__zz_regVec_0 = regVec_3326;
      end
      12'b110011111111 : begin
        _zz__zz_regVec_0 = regVec_3327;
      end
      12'b110100000000 : begin
        _zz__zz_regVec_0 = regVec_3328;
      end
      12'b110100000001 : begin
        _zz__zz_regVec_0 = regVec_3329;
      end
      12'b110100000010 : begin
        _zz__zz_regVec_0 = regVec_3330;
      end
      12'b110100000011 : begin
        _zz__zz_regVec_0 = regVec_3331;
      end
      12'b110100000100 : begin
        _zz__zz_regVec_0 = regVec_3332;
      end
      12'b110100000101 : begin
        _zz__zz_regVec_0 = regVec_3333;
      end
      12'b110100000110 : begin
        _zz__zz_regVec_0 = regVec_3334;
      end
      12'b110100000111 : begin
        _zz__zz_regVec_0 = regVec_3335;
      end
      12'b110100001000 : begin
        _zz__zz_regVec_0 = regVec_3336;
      end
      12'b110100001001 : begin
        _zz__zz_regVec_0 = regVec_3337;
      end
      12'b110100001010 : begin
        _zz__zz_regVec_0 = regVec_3338;
      end
      12'b110100001011 : begin
        _zz__zz_regVec_0 = regVec_3339;
      end
      12'b110100001100 : begin
        _zz__zz_regVec_0 = regVec_3340;
      end
      12'b110100001101 : begin
        _zz__zz_regVec_0 = regVec_3341;
      end
      12'b110100001110 : begin
        _zz__zz_regVec_0 = regVec_3342;
      end
      12'b110100001111 : begin
        _zz__zz_regVec_0 = regVec_3343;
      end
      12'b110100010000 : begin
        _zz__zz_regVec_0 = regVec_3344;
      end
      12'b110100010001 : begin
        _zz__zz_regVec_0 = regVec_3345;
      end
      12'b110100010010 : begin
        _zz__zz_regVec_0 = regVec_3346;
      end
      12'b110100010011 : begin
        _zz__zz_regVec_0 = regVec_3347;
      end
      12'b110100010100 : begin
        _zz__zz_regVec_0 = regVec_3348;
      end
      12'b110100010101 : begin
        _zz__zz_regVec_0 = regVec_3349;
      end
      12'b110100010110 : begin
        _zz__zz_regVec_0 = regVec_3350;
      end
      12'b110100010111 : begin
        _zz__zz_regVec_0 = regVec_3351;
      end
      12'b110100011000 : begin
        _zz__zz_regVec_0 = regVec_3352;
      end
      12'b110100011001 : begin
        _zz__zz_regVec_0 = regVec_3353;
      end
      12'b110100011010 : begin
        _zz__zz_regVec_0 = regVec_3354;
      end
      12'b110100011011 : begin
        _zz__zz_regVec_0 = regVec_3355;
      end
      12'b110100011100 : begin
        _zz__zz_regVec_0 = regVec_3356;
      end
      12'b110100011101 : begin
        _zz__zz_regVec_0 = regVec_3357;
      end
      12'b110100011110 : begin
        _zz__zz_regVec_0 = regVec_3358;
      end
      12'b110100011111 : begin
        _zz__zz_regVec_0 = regVec_3359;
      end
      12'b110100100000 : begin
        _zz__zz_regVec_0 = regVec_3360;
      end
      12'b110100100001 : begin
        _zz__zz_regVec_0 = regVec_3361;
      end
      12'b110100100010 : begin
        _zz__zz_regVec_0 = regVec_3362;
      end
      12'b110100100011 : begin
        _zz__zz_regVec_0 = regVec_3363;
      end
      12'b110100100100 : begin
        _zz__zz_regVec_0 = regVec_3364;
      end
      12'b110100100101 : begin
        _zz__zz_regVec_0 = regVec_3365;
      end
      12'b110100100110 : begin
        _zz__zz_regVec_0 = regVec_3366;
      end
      12'b110100100111 : begin
        _zz__zz_regVec_0 = regVec_3367;
      end
      12'b110100101000 : begin
        _zz__zz_regVec_0 = regVec_3368;
      end
      12'b110100101001 : begin
        _zz__zz_regVec_0 = regVec_3369;
      end
      12'b110100101010 : begin
        _zz__zz_regVec_0 = regVec_3370;
      end
      12'b110100101011 : begin
        _zz__zz_regVec_0 = regVec_3371;
      end
      12'b110100101100 : begin
        _zz__zz_regVec_0 = regVec_3372;
      end
      12'b110100101101 : begin
        _zz__zz_regVec_0 = regVec_3373;
      end
      12'b110100101110 : begin
        _zz__zz_regVec_0 = regVec_3374;
      end
      12'b110100101111 : begin
        _zz__zz_regVec_0 = regVec_3375;
      end
      12'b110100110000 : begin
        _zz__zz_regVec_0 = regVec_3376;
      end
      12'b110100110001 : begin
        _zz__zz_regVec_0 = regVec_3377;
      end
      12'b110100110010 : begin
        _zz__zz_regVec_0 = regVec_3378;
      end
      12'b110100110011 : begin
        _zz__zz_regVec_0 = regVec_3379;
      end
      12'b110100110100 : begin
        _zz__zz_regVec_0 = regVec_3380;
      end
      12'b110100110101 : begin
        _zz__zz_regVec_0 = regVec_3381;
      end
      12'b110100110110 : begin
        _zz__zz_regVec_0 = regVec_3382;
      end
      12'b110100110111 : begin
        _zz__zz_regVec_0 = regVec_3383;
      end
      12'b110100111000 : begin
        _zz__zz_regVec_0 = regVec_3384;
      end
      12'b110100111001 : begin
        _zz__zz_regVec_0 = regVec_3385;
      end
      12'b110100111010 : begin
        _zz__zz_regVec_0 = regVec_3386;
      end
      12'b110100111011 : begin
        _zz__zz_regVec_0 = regVec_3387;
      end
      12'b110100111100 : begin
        _zz__zz_regVec_0 = regVec_3388;
      end
      12'b110100111101 : begin
        _zz__zz_regVec_0 = regVec_3389;
      end
      12'b110100111110 : begin
        _zz__zz_regVec_0 = regVec_3390;
      end
      12'b110100111111 : begin
        _zz__zz_regVec_0 = regVec_3391;
      end
      12'b110101000000 : begin
        _zz__zz_regVec_0 = regVec_3392;
      end
      12'b110101000001 : begin
        _zz__zz_regVec_0 = regVec_3393;
      end
      12'b110101000010 : begin
        _zz__zz_regVec_0 = regVec_3394;
      end
      12'b110101000011 : begin
        _zz__zz_regVec_0 = regVec_3395;
      end
      12'b110101000100 : begin
        _zz__zz_regVec_0 = regVec_3396;
      end
      12'b110101000101 : begin
        _zz__zz_regVec_0 = regVec_3397;
      end
      12'b110101000110 : begin
        _zz__zz_regVec_0 = regVec_3398;
      end
      12'b110101000111 : begin
        _zz__zz_regVec_0 = regVec_3399;
      end
      12'b110101001000 : begin
        _zz__zz_regVec_0 = regVec_3400;
      end
      12'b110101001001 : begin
        _zz__zz_regVec_0 = regVec_3401;
      end
      12'b110101001010 : begin
        _zz__zz_regVec_0 = regVec_3402;
      end
      12'b110101001011 : begin
        _zz__zz_regVec_0 = regVec_3403;
      end
      12'b110101001100 : begin
        _zz__zz_regVec_0 = regVec_3404;
      end
      12'b110101001101 : begin
        _zz__zz_regVec_0 = regVec_3405;
      end
      12'b110101001110 : begin
        _zz__zz_regVec_0 = regVec_3406;
      end
      12'b110101001111 : begin
        _zz__zz_regVec_0 = regVec_3407;
      end
      12'b110101010000 : begin
        _zz__zz_regVec_0 = regVec_3408;
      end
      12'b110101010001 : begin
        _zz__zz_regVec_0 = regVec_3409;
      end
      12'b110101010010 : begin
        _zz__zz_regVec_0 = regVec_3410;
      end
      12'b110101010011 : begin
        _zz__zz_regVec_0 = regVec_3411;
      end
      12'b110101010100 : begin
        _zz__zz_regVec_0 = regVec_3412;
      end
      12'b110101010101 : begin
        _zz__zz_regVec_0 = regVec_3413;
      end
      12'b110101010110 : begin
        _zz__zz_regVec_0 = regVec_3414;
      end
      12'b110101010111 : begin
        _zz__zz_regVec_0 = regVec_3415;
      end
      12'b110101011000 : begin
        _zz__zz_regVec_0 = regVec_3416;
      end
      12'b110101011001 : begin
        _zz__zz_regVec_0 = regVec_3417;
      end
      12'b110101011010 : begin
        _zz__zz_regVec_0 = regVec_3418;
      end
      12'b110101011011 : begin
        _zz__zz_regVec_0 = regVec_3419;
      end
      12'b110101011100 : begin
        _zz__zz_regVec_0 = regVec_3420;
      end
      12'b110101011101 : begin
        _zz__zz_regVec_0 = regVec_3421;
      end
      12'b110101011110 : begin
        _zz__zz_regVec_0 = regVec_3422;
      end
      12'b110101011111 : begin
        _zz__zz_regVec_0 = regVec_3423;
      end
      12'b110101100000 : begin
        _zz__zz_regVec_0 = regVec_3424;
      end
      12'b110101100001 : begin
        _zz__zz_regVec_0 = regVec_3425;
      end
      12'b110101100010 : begin
        _zz__zz_regVec_0 = regVec_3426;
      end
      12'b110101100011 : begin
        _zz__zz_regVec_0 = regVec_3427;
      end
      12'b110101100100 : begin
        _zz__zz_regVec_0 = regVec_3428;
      end
      12'b110101100101 : begin
        _zz__zz_regVec_0 = regVec_3429;
      end
      12'b110101100110 : begin
        _zz__zz_regVec_0 = regVec_3430;
      end
      12'b110101100111 : begin
        _zz__zz_regVec_0 = regVec_3431;
      end
      12'b110101101000 : begin
        _zz__zz_regVec_0 = regVec_3432;
      end
      12'b110101101001 : begin
        _zz__zz_regVec_0 = regVec_3433;
      end
      12'b110101101010 : begin
        _zz__zz_regVec_0 = regVec_3434;
      end
      12'b110101101011 : begin
        _zz__zz_regVec_0 = regVec_3435;
      end
      12'b110101101100 : begin
        _zz__zz_regVec_0 = regVec_3436;
      end
      12'b110101101101 : begin
        _zz__zz_regVec_0 = regVec_3437;
      end
      12'b110101101110 : begin
        _zz__zz_regVec_0 = regVec_3438;
      end
      12'b110101101111 : begin
        _zz__zz_regVec_0 = regVec_3439;
      end
      12'b110101110000 : begin
        _zz__zz_regVec_0 = regVec_3440;
      end
      12'b110101110001 : begin
        _zz__zz_regVec_0 = regVec_3441;
      end
      12'b110101110010 : begin
        _zz__zz_regVec_0 = regVec_3442;
      end
      12'b110101110011 : begin
        _zz__zz_regVec_0 = regVec_3443;
      end
      12'b110101110100 : begin
        _zz__zz_regVec_0 = regVec_3444;
      end
      12'b110101110101 : begin
        _zz__zz_regVec_0 = regVec_3445;
      end
      12'b110101110110 : begin
        _zz__zz_regVec_0 = regVec_3446;
      end
      12'b110101110111 : begin
        _zz__zz_regVec_0 = regVec_3447;
      end
      12'b110101111000 : begin
        _zz__zz_regVec_0 = regVec_3448;
      end
      12'b110101111001 : begin
        _zz__zz_regVec_0 = regVec_3449;
      end
      12'b110101111010 : begin
        _zz__zz_regVec_0 = regVec_3450;
      end
      12'b110101111011 : begin
        _zz__zz_regVec_0 = regVec_3451;
      end
      12'b110101111100 : begin
        _zz__zz_regVec_0 = regVec_3452;
      end
      12'b110101111101 : begin
        _zz__zz_regVec_0 = regVec_3453;
      end
      12'b110101111110 : begin
        _zz__zz_regVec_0 = regVec_3454;
      end
      12'b110101111111 : begin
        _zz__zz_regVec_0 = regVec_3455;
      end
      12'b110110000000 : begin
        _zz__zz_regVec_0 = regVec_3456;
      end
      12'b110110000001 : begin
        _zz__zz_regVec_0 = regVec_3457;
      end
      12'b110110000010 : begin
        _zz__zz_regVec_0 = regVec_3458;
      end
      12'b110110000011 : begin
        _zz__zz_regVec_0 = regVec_3459;
      end
      12'b110110000100 : begin
        _zz__zz_regVec_0 = regVec_3460;
      end
      12'b110110000101 : begin
        _zz__zz_regVec_0 = regVec_3461;
      end
      12'b110110000110 : begin
        _zz__zz_regVec_0 = regVec_3462;
      end
      12'b110110000111 : begin
        _zz__zz_regVec_0 = regVec_3463;
      end
      12'b110110001000 : begin
        _zz__zz_regVec_0 = regVec_3464;
      end
      12'b110110001001 : begin
        _zz__zz_regVec_0 = regVec_3465;
      end
      12'b110110001010 : begin
        _zz__zz_regVec_0 = regVec_3466;
      end
      12'b110110001011 : begin
        _zz__zz_regVec_0 = regVec_3467;
      end
      12'b110110001100 : begin
        _zz__zz_regVec_0 = regVec_3468;
      end
      12'b110110001101 : begin
        _zz__zz_regVec_0 = regVec_3469;
      end
      12'b110110001110 : begin
        _zz__zz_regVec_0 = regVec_3470;
      end
      12'b110110001111 : begin
        _zz__zz_regVec_0 = regVec_3471;
      end
      12'b110110010000 : begin
        _zz__zz_regVec_0 = regVec_3472;
      end
      12'b110110010001 : begin
        _zz__zz_regVec_0 = regVec_3473;
      end
      12'b110110010010 : begin
        _zz__zz_regVec_0 = regVec_3474;
      end
      12'b110110010011 : begin
        _zz__zz_regVec_0 = regVec_3475;
      end
      12'b110110010100 : begin
        _zz__zz_regVec_0 = regVec_3476;
      end
      12'b110110010101 : begin
        _zz__zz_regVec_0 = regVec_3477;
      end
      12'b110110010110 : begin
        _zz__zz_regVec_0 = regVec_3478;
      end
      12'b110110010111 : begin
        _zz__zz_regVec_0 = regVec_3479;
      end
      12'b110110011000 : begin
        _zz__zz_regVec_0 = regVec_3480;
      end
      12'b110110011001 : begin
        _zz__zz_regVec_0 = regVec_3481;
      end
      12'b110110011010 : begin
        _zz__zz_regVec_0 = regVec_3482;
      end
      12'b110110011011 : begin
        _zz__zz_regVec_0 = regVec_3483;
      end
      12'b110110011100 : begin
        _zz__zz_regVec_0 = regVec_3484;
      end
      12'b110110011101 : begin
        _zz__zz_regVec_0 = regVec_3485;
      end
      12'b110110011110 : begin
        _zz__zz_regVec_0 = regVec_3486;
      end
      12'b110110011111 : begin
        _zz__zz_regVec_0 = regVec_3487;
      end
      12'b110110100000 : begin
        _zz__zz_regVec_0 = regVec_3488;
      end
      12'b110110100001 : begin
        _zz__zz_regVec_0 = regVec_3489;
      end
      12'b110110100010 : begin
        _zz__zz_regVec_0 = regVec_3490;
      end
      12'b110110100011 : begin
        _zz__zz_regVec_0 = regVec_3491;
      end
      12'b110110100100 : begin
        _zz__zz_regVec_0 = regVec_3492;
      end
      12'b110110100101 : begin
        _zz__zz_regVec_0 = regVec_3493;
      end
      12'b110110100110 : begin
        _zz__zz_regVec_0 = regVec_3494;
      end
      12'b110110100111 : begin
        _zz__zz_regVec_0 = regVec_3495;
      end
      12'b110110101000 : begin
        _zz__zz_regVec_0 = regVec_3496;
      end
      12'b110110101001 : begin
        _zz__zz_regVec_0 = regVec_3497;
      end
      12'b110110101010 : begin
        _zz__zz_regVec_0 = regVec_3498;
      end
      12'b110110101011 : begin
        _zz__zz_regVec_0 = regVec_3499;
      end
      12'b110110101100 : begin
        _zz__zz_regVec_0 = regVec_3500;
      end
      12'b110110101101 : begin
        _zz__zz_regVec_0 = regVec_3501;
      end
      12'b110110101110 : begin
        _zz__zz_regVec_0 = regVec_3502;
      end
      12'b110110101111 : begin
        _zz__zz_regVec_0 = regVec_3503;
      end
      12'b110110110000 : begin
        _zz__zz_regVec_0 = regVec_3504;
      end
      12'b110110110001 : begin
        _zz__zz_regVec_0 = regVec_3505;
      end
      12'b110110110010 : begin
        _zz__zz_regVec_0 = regVec_3506;
      end
      12'b110110110011 : begin
        _zz__zz_regVec_0 = regVec_3507;
      end
      12'b110110110100 : begin
        _zz__zz_regVec_0 = regVec_3508;
      end
      12'b110110110101 : begin
        _zz__zz_regVec_0 = regVec_3509;
      end
      12'b110110110110 : begin
        _zz__zz_regVec_0 = regVec_3510;
      end
      12'b110110110111 : begin
        _zz__zz_regVec_0 = regVec_3511;
      end
      12'b110110111000 : begin
        _zz__zz_regVec_0 = regVec_3512;
      end
      12'b110110111001 : begin
        _zz__zz_regVec_0 = regVec_3513;
      end
      12'b110110111010 : begin
        _zz__zz_regVec_0 = regVec_3514;
      end
      12'b110110111011 : begin
        _zz__zz_regVec_0 = regVec_3515;
      end
      12'b110110111100 : begin
        _zz__zz_regVec_0 = regVec_3516;
      end
      12'b110110111101 : begin
        _zz__zz_regVec_0 = regVec_3517;
      end
      12'b110110111110 : begin
        _zz__zz_regVec_0 = regVec_3518;
      end
      12'b110110111111 : begin
        _zz__zz_regVec_0 = regVec_3519;
      end
      12'b110111000000 : begin
        _zz__zz_regVec_0 = regVec_3520;
      end
      12'b110111000001 : begin
        _zz__zz_regVec_0 = regVec_3521;
      end
      12'b110111000010 : begin
        _zz__zz_regVec_0 = regVec_3522;
      end
      12'b110111000011 : begin
        _zz__zz_regVec_0 = regVec_3523;
      end
      12'b110111000100 : begin
        _zz__zz_regVec_0 = regVec_3524;
      end
      12'b110111000101 : begin
        _zz__zz_regVec_0 = regVec_3525;
      end
      12'b110111000110 : begin
        _zz__zz_regVec_0 = regVec_3526;
      end
      12'b110111000111 : begin
        _zz__zz_regVec_0 = regVec_3527;
      end
      12'b110111001000 : begin
        _zz__zz_regVec_0 = regVec_3528;
      end
      12'b110111001001 : begin
        _zz__zz_regVec_0 = regVec_3529;
      end
      12'b110111001010 : begin
        _zz__zz_regVec_0 = regVec_3530;
      end
      12'b110111001011 : begin
        _zz__zz_regVec_0 = regVec_3531;
      end
      12'b110111001100 : begin
        _zz__zz_regVec_0 = regVec_3532;
      end
      12'b110111001101 : begin
        _zz__zz_regVec_0 = regVec_3533;
      end
      12'b110111001110 : begin
        _zz__zz_regVec_0 = regVec_3534;
      end
      12'b110111001111 : begin
        _zz__zz_regVec_0 = regVec_3535;
      end
      12'b110111010000 : begin
        _zz__zz_regVec_0 = regVec_3536;
      end
      12'b110111010001 : begin
        _zz__zz_regVec_0 = regVec_3537;
      end
      12'b110111010010 : begin
        _zz__zz_regVec_0 = regVec_3538;
      end
      12'b110111010011 : begin
        _zz__zz_regVec_0 = regVec_3539;
      end
      12'b110111010100 : begin
        _zz__zz_regVec_0 = regVec_3540;
      end
      12'b110111010101 : begin
        _zz__zz_regVec_0 = regVec_3541;
      end
      12'b110111010110 : begin
        _zz__zz_regVec_0 = regVec_3542;
      end
      12'b110111010111 : begin
        _zz__zz_regVec_0 = regVec_3543;
      end
      12'b110111011000 : begin
        _zz__zz_regVec_0 = regVec_3544;
      end
      12'b110111011001 : begin
        _zz__zz_regVec_0 = regVec_3545;
      end
      12'b110111011010 : begin
        _zz__zz_regVec_0 = regVec_3546;
      end
      12'b110111011011 : begin
        _zz__zz_regVec_0 = regVec_3547;
      end
      12'b110111011100 : begin
        _zz__zz_regVec_0 = regVec_3548;
      end
      12'b110111011101 : begin
        _zz__zz_regVec_0 = regVec_3549;
      end
      12'b110111011110 : begin
        _zz__zz_regVec_0 = regVec_3550;
      end
      12'b110111011111 : begin
        _zz__zz_regVec_0 = regVec_3551;
      end
      12'b110111100000 : begin
        _zz__zz_regVec_0 = regVec_3552;
      end
      12'b110111100001 : begin
        _zz__zz_regVec_0 = regVec_3553;
      end
      12'b110111100010 : begin
        _zz__zz_regVec_0 = regVec_3554;
      end
      12'b110111100011 : begin
        _zz__zz_regVec_0 = regVec_3555;
      end
      12'b110111100100 : begin
        _zz__zz_regVec_0 = regVec_3556;
      end
      12'b110111100101 : begin
        _zz__zz_regVec_0 = regVec_3557;
      end
      12'b110111100110 : begin
        _zz__zz_regVec_0 = regVec_3558;
      end
      12'b110111100111 : begin
        _zz__zz_regVec_0 = regVec_3559;
      end
      12'b110111101000 : begin
        _zz__zz_regVec_0 = regVec_3560;
      end
      12'b110111101001 : begin
        _zz__zz_regVec_0 = regVec_3561;
      end
      12'b110111101010 : begin
        _zz__zz_regVec_0 = regVec_3562;
      end
      12'b110111101011 : begin
        _zz__zz_regVec_0 = regVec_3563;
      end
      12'b110111101100 : begin
        _zz__zz_regVec_0 = regVec_3564;
      end
      12'b110111101101 : begin
        _zz__zz_regVec_0 = regVec_3565;
      end
      12'b110111101110 : begin
        _zz__zz_regVec_0 = regVec_3566;
      end
      12'b110111101111 : begin
        _zz__zz_regVec_0 = regVec_3567;
      end
      12'b110111110000 : begin
        _zz__zz_regVec_0 = regVec_3568;
      end
      12'b110111110001 : begin
        _zz__zz_regVec_0 = regVec_3569;
      end
      12'b110111110010 : begin
        _zz__zz_regVec_0 = regVec_3570;
      end
      12'b110111110011 : begin
        _zz__zz_regVec_0 = regVec_3571;
      end
      12'b110111110100 : begin
        _zz__zz_regVec_0 = regVec_3572;
      end
      12'b110111110101 : begin
        _zz__zz_regVec_0 = regVec_3573;
      end
      12'b110111110110 : begin
        _zz__zz_regVec_0 = regVec_3574;
      end
      12'b110111110111 : begin
        _zz__zz_regVec_0 = regVec_3575;
      end
      12'b110111111000 : begin
        _zz__zz_regVec_0 = regVec_3576;
      end
      12'b110111111001 : begin
        _zz__zz_regVec_0 = regVec_3577;
      end
      12'b110111111010 : begin
        _zz__zz_regVec_0 = regVec_3578;
      end
      12'b110111111011 : begin
        _zz__zz_regVec_0 = regVec_3579;
      end
      12'b110111111100 : begin
        _zz__zz_regVec_0 = regVec_3580;
      end
      12'b110111111101 : begin
        _zz__zz_regVec_0 = regVec_3581;
      end
      12'b110111111110 : begin
        _zz__zz_regVec_0 = regVec_3582;
      end
      12'b110111111111 : begin
        _zz__zz_regVec_0 = regVec_3583;
      end
      12'b111000000000 : begin
        _zz__zz_regVec_0 = regVec_3584;
      end
      12'b111000000001 : begin
        _zz__zz_regVec_0 = regVec_3585;
      end
      12'b111000000010 : begin
        _zz__zz_regVec_0 = regVec_3586;
      end
      12'b111000000011 : begin
        _zz__zz_regVec_0 = regVec_3587;
      end
      12'b111000000100 : begin
        _zz__zz_regVec_0 = regVec_3588;
      end
      12'b111000000101 : begin
        _zz__zz_regVec_0 = regVec_3589;
      end
      12'b111000000110 : begin
        _zz__zz_regVec_0 = regVec_3590;
      end
      12'b111000000111 : begin
        _zz__zz_regVec_0 = regVec_3591;
      end
      12'b111000001000 : begin
        _zz__zz_regVec_0 = regVec_3592;
      end
      12'b111000001001 : begin
        _zz__zz_regVec_0 = regVec_3593;
      end
      12'b111000001010 : begin
        _zz__zz_regVec_0 = regVec_3594;
      end
      12'b111000001011 : begin
        _zz__zz_regVec_0 = regVec_3595;
      end
      12'b111000001100 : begin
        _zz__zz_regVec_0 = regVec_3596;
      end
      12'b111000001101 : begin
        _zz__zz_regVec_0 = regVec_3597;
      end
      12'b111000001110 : begin
        _zz__zz_regVec_0 = regVec_3598;
      end
      12'b111000001111 : begin
        _zz__zz_regVec_0 = regVec_3599;
      end
      12'b111000010000 : begin
        _zz__zz_regVec_0 = regVec_3600;
      end
      12'b111000010001 : begin
        _zz__zz_regVec_0 = regVec_3601;
      end
      12'b111000010010 : begin
        _zz__zz_regVec_0 = regVec_3602;
      end
      12'b111000010011 : begin
        _zz__zz_regVec_0 = regVec_3603;
      end
      12'b111000010100 : begin
        _zz__zz_regVec_0 = regVec_3604;
      end
      12'b111000010101 : begin
        _zz__zz_regVec_0 = regVec_3605;
      end
      12'b111000010110 : begin
        _zz__zz_regVec_0 = regVec_3606;
      end
      12'b111000010111 : begin
        _zz__zz_regVec_0 = regVec_3607;
      end
      12'b111000011000 : begin
        _zz__zz_regVec_0 = regVec_3608;
      end
      12'b111000011001 : begin
        _zz__zz_regVec_0 = regVec_3609;
      end
      12'b111000011010 : begin
        _zz__zz_regVec_0 = regVec_3610;
      end
      12'b111000011011 : begin
        _zz__zz_regVec_0 = regVec_3611;
      end
      12'b111000011100 : begin
        _zz__zz_regVec_0 = regVec_3612;
      end
      12'b111000011101 : begin
        _zz__zz_regVec_0 = regVec_3613;
      end
      12'b111000011110 : begin
        _zz__zz_regVec_0 = regVec_3614;
      end
      12'b111000011111 : begin
        _zz__zz_regVec_0 = regVec_3615;
      end
      12'b111000100000 : begin
        _zz__zz_regVec_0 = regVec_3616;
      end
      12'b111000100001 : begin
        _zz__zz_regVec_0 = regVec_3617;
      end
      12'b111000100010 : begin
        _zz__zz_regVec_0 = regVec_3618;
      end
      12'b111000100011 : begin
        _zz__zz_regVec_0 = regVec_3619;
      end
      12'b111000100100 : begin
        _zz__zz_regVec_0 = regVec_3620;
      end
      12'b111000100101 : begin
        _zz__zz_regVec_0 = regVec_3621;
      end
      12'b111000100110 : begin
        _zz__zz_regVec_0 = regVec_3622;
      end
      12'b111000100111 : begin
        _zz__zz_regVec_0 = regVec_3623;
      end
      12'b111000101000 : begin
        _zz__zz_regVec_0 = regVec_3624;
      end
      12'b111000101001 : begin
        _zz__zz_regVec_0 = regVec_3625;
      end
      12'b111000101010 : begin
        _zz__zz_regVec_0 = regVec_3626;
      end
      12'b111000101011 : begin
        _zz__zz_regVec_0 = regVec_3627;
      end
      12'b111000101100 : begin
        _zz__zz_regVec_0 = regVec_3628;
      end
      12'b111000101101 : begin
        _zz__zz_regVec_0 = regVec_3629;
      end
      12'b111000101110 : begin
        _zz__zz_regVec_0 = regVec_3630;
      end
      12'b111000101111 : begin
        _zz__zz_regVec_0 = regVec_3631;
      end
      12'b111000110000 : begin
        _zz__zz_regVec_0 = regVec_3632;
      end
      12'b111000110001 : begin
        _zz__zz_regVec_0 = regVec_3633;
      end
      12'b111000110010 : begin
        _zz__zz_regVec_0 = regVec_3634;
      end
      12'b111000110011 : begin
        _zz__zz_regVec_0 = regVec_3635;
      end
      12'b111000110100 : begin
        _zz__zz_regVec_0 = regVec_3636;
      end
      12'b111000110101 : begin
        _zz__zz_regVec_0 = regVec_3637;
      end
      12'b111000110110 : begin
        _zz__zz_regVec_0 = regVec_3638;
      end
      12'b111000110111 : begin
        _zz__zz_regVec_0 = regVec_3639;
      end
      12'b111000111000 : begin
        _zz__zz_regVec_0 = regVec_3640;
      end
      12'b111000111001 : begin
        _zz__zz_regVec_0 = regVec_3641;
      end
      12'b111000111010 : begin
        _zz__zz_regVec_0 = regVec_3642;
      end
      12'b111000111011 : begin
        _zz__zz_regVec_0 = regVec_3643;
      end
      12'b111000111100 : begin
        _zz__zz_regVec_0 = regVec_3644;
      end
      12'b111000111101 : begin
        _zz__zz_regVec_0 = regVec_3645;
      end
      12'b111000111110 : begin
        _zz__zz_regVec_0 = regVec_3646;
      end
      12'b111000111111 : begin
        _zz__zz_regVec_0 = regVec_3647;
      end
      12'b111001000000 : begin
        _zz__zz_regVec_0 = regVec_3648;
      end
      12'b111001000001 : begin
        _zz__zz_regVec_0 = regVec_3649;
      end
      12'b111001000010 : begin
        _zz__zz_regVec_0 = regVec_3650;
      end
      12'b111001000011 : begin
        _zz__zz_regVec_0 = regVec_3651;
      end
      12'b111001000100 : begin
        _zz__zz_regVec_0 = regVec_3652;
      end
      12'b111001000101 : begin
        _zz__zz_regVec_0 = regVec_3653;
      end
      12'b111001000110 : begin
        _zz__zz_regVec_0 = regVec_3654;
      end
      12'b111001000111 : begin
        _zz__zz_regVec_0 = regVec_3655;
      end
      12'b111001001000 : begin
        _zz__zz_regVec_0 = regVec_3656;
      end
      12'b111001001001 : begin
        _zz__zz_regVec_0 = regVec_3657;
      end
      12'b111001001010 : begin
        _zz__zz_regVec_0 = regVec_3658;
      end
      12'b111001001011 : begin
        _zz__zz_regVec_0 = regVec_3659;
      end
      12'b111001001100 : begin
        _zz__zz_regVec_0 = regVec_3660;
      end
      12'b111001001101 : begin
        _zz__zz_regVec_0 = regVec_3661;
      end
      12'b111001001110 : begin
        _zz__zz_regVec_0 = regVec_3662;
      end
      12'b111001001111 : begin
        _zz__zz_regVec_0 = regVec_3663;
      end
      12'b111001010000 : begin
        _zz__zz_regVec_0 = regVec_3664;
      end
      12'b111001010001 : begin
        _zz__zz_regVec_0 = regVec_3665;
      end
      12'b111001010010 : begin
        _zz__zz_regVec_0 = regVec_3666;
      end
      12'b111001010011 : begin
        _zz__zz_regVec_0 = regVec_3667;
      end
      12'b111001010100 : begin
        _zz__zz_regVec_0 = regVec_3668;
      end
      12'b111001010101 : begin
        _zz__zz_regVec_0 = regVec_3669;
      end
      12'b111001010110 : begin
        _zz__zz_regVec_0 = regVec_3670;
      end
      12'b111001010111 : begin
        _zz__zz_regVec_0 = regVec_3671;
      end
      12'b111001011000 : begin
        _zz__zz_regVec_0 = regVec_3672;
      end
      12'b111001011001 : begin
        _zz__zz_regVec_0 = regVec_3673;
      end
      12'b111001011010 : begin
        _zz__zz_regVec_0 = regVec_3674;
      end
      12'b111001011011 : begin
        _zz__zz_regVec_0 = regVec_3675;
      end
      12'b111001011100 : begin
        _zz__zz_regVec_0 = regVec_3676;
      end
      12'b111001011101 : begin
        _zz__zz_regVec_0 = regVec_3677;
      end
      12'b111001011110 : begin
        _zz__zz_regVec_0 = regVec_3678;
      end
      12'b111001011111 : begin
        _zz__zz_regVec_0 = regVec_3679;
      end
      12'b111001100000 : begin
        _zz__zz_regVec_0 = regVec_3680;
      end
      12'b111001100001 : begin
        _zz__zz_regVec_0 = regVec_3681;
      end
      12'b111001100010 : begin
        _zz__zz_regVec_0 = regVec_3682;
      end
      12'b111001100011 : begin
        _zz__zz_regVec_0 = regVec_3683;
      end
      12'b111001100100 : begin
        _zz__zz_regVec_0 = regVec_3684;
      end
      12'b111001100101 : begin
        _zz__zz_regVec_0 = regVec_3685;
      end
      12'b111001100110 : begin
        _zz__zz_regVec_0 = regVec_3686;
      end
      12'b111001100111 : begin
        _zz__zz_regVec_0 = regVec_3687;
      end
      12'b111001101000 : begin
        _zz__zz_regVec_0 = regVec_3688;
      end
      12'b111001101001 : begin
        _zz__zz_regVec_0 = regVec_3689;
      end
      12'b111001101010 : begin
        _zz__zz_regVec_0 = regVec_3690;
      end
      12'b111001101011 : begin
        _zz__zz_regVec_0 = regVec_3691;
      end
      12'b111001101100 : begin
        _zz__zz_regVec_0 = regVec_3692;
      end
      12'b111001101101 : begin
        _zz__zz_regVec_0 = regVec_3693;
      end
      12'b111001101110 : begin
        _zz__zz_regVec_0 = regVec_3694;
      end
      12'b111001101111 : begin
        _zz__zz_regVec_0 = regVec_3695;
      end
      12'b111001110000 : begin
        _zz__zz_regVec_0 = regVec_3696;
      end
      12'b111001110001 : begin
        _zz__zz_regVec_0 = regVec_3697;
      end
      12'b111001110010 : begin
        _zz__zz_regVec_0 = regVec_3698;
      end
      12'b111001110011 : begin
        _zz__zz_regVec_0 = regVec_3699;
      end
      12'b111001110100 : begin
        _zz__zz_regVec_0 = regVec_3700;
      end
      12'b111001110101 : begin
        _zz__zz_regVec_0 = regVec_3701;
      end
      12'b111001110110 : begin
        _zz__zz_regVec_0 = regVec_3702;
      end
      12'b111001110111 : begin
        _zz__zz_regVec_0 = regVec_3703;
      end
      12'b111001111000 : begin
        _zz__zz_regVec_0 = regVec_3704;
      end
      12'b111001111001 : begin
        _zz__zz_regVec_0 = regVec_3705;
      end
      12'b111001111010 : begin
        _zz__zz_regVec_0 = regVec_3706;
      end
      12'b111001111011 : begin
        _zz__zz_regVec_0 = regVec_3707;
      end
      12'b111001111100 : begin
        _zz__zz_regVec_0 = regVec_3708;
      end
      12'b111001111101 : begin
        _zz__zz_regVec_0 = regVec_3709;
      end
      12'b111001111110 : begin
        _zz__zz_regVec_0 = regVec_3710;
      end
      12'b111001111111 : begin
        _zz__zz_regVec_0 = regVec_3711;
      end
      12'b111010000000 : begin
        _zz__zz_regVec_0 = regVec_3712;
      end
      12'b111010000001 : begin
        _zz__zz_regVec_0 = regVec_3713;
      end
      12'b111010000010 : begin
        _zz__zz_regVec_0 = regVec_3714;
      end
      12'b111010000011 : begin
        _zz__zz_regVec_0 = regVec_3715;
      end
      12'b111010000100 : begin
        _zz__zz_regVec_0 = regVec_3716;
      end
      12'b111010000101 : begin
        _zz__zz_regVec_0 = regVec_3717;
      end
      12'b111010000110 : begin
        _zz__zz_regVec_0 = regVec_3718;
      end
      12'b111010000111 : begin
        _zz__zz_regVec_0 = regVec_3719;
      end
      12'b111010001000 : begin
        _zz__zz_regVec_0 = regVec_3720;
      end
      12'b111010001001 : begin
        _zz__zz_regVec_0 = regVec_3721;
      end
      12'b111010001010 : begin
        _zz__zz_regVec_0 = regVec_3722;
      end
      12'b111010001011 : begin
        _zz__zz_regVec_0 = regVec_3723;
      end
      12'b111010001100 : begin
        _zz__zz_regVec_0 = regVec_3724;
      end
      12'b111010001101 : begin
        _zz__zz_regVec_0 = regVec_3725;
      end
      12'b111010001110 : begin
        _zz__zz_regVec_0 = regVec_3726;
      end
      12'b111010001111 : begin
        _zz__zz_regVec_0 = regVec_3727;
      end
      12'b111010010000 : begin
        _zz__zz_regVec_0 = regVec_3728;
      end
      12'b111010010001 : begin
        _zz__zz_regVec_0 = regVec_3729;
      end
      12'b111010010010 : begin
        _zz__zz_regVec_0 = regVec_3730;
      end
      12'b111010010011 : begin
        _zz__zz_regVec_0 = regVec_3731;
      end
      12'b111010010100 : begin
        _zz__zz_regVec_0 = regVec_3732;
      end
      12'b111010010101 : begin
        _zz__zz_regVec_0 = regVec_3733;
      end
      12'b111010010110 : begin
        _zz__zz_regVec_0 = regVec_3734;
      end
      12'b111010010111 : begin
        _zz__zz_regVec_0 = regVec_3735;
      end
      12'b111010011000 : begin
        _zz__zz_regVec_0 = regVec_3736;
      end
      12'b111010011001 : begin
        _zz__zz_regVec_0 = regVec_3737;
      end
      12'b111010011010 : begin
        _zz__zz_regVec_0 = regVec_3738;
      end
      12'b111010011011 : begin
        _zz__zz_regVec_0 = regVec_3739;
      end
      12'b111010011100 : begin
        _zz__zz_regVec_0 = regVec_3740;
      end
      12'b111010011101 : begin
        _zz__zz_regVec_0 = regVec_3741;
      end
      12'b111010011110 : begin
        _zz__zz_regVec_0 = regVec_3742;
      end
      12'b111010011111 : begin
        _zz__zz_regVec_0 = regVec_3743;
      end
      12'b111010100000 : begin
        _zz__zz_regVec_0 = regVec_3744;
      end
      12'b111010100001 : begin
        _zz__zz_regVec_0 = regVec_3745;
      end
      12'b111010100010 : begin
        _zz__zz_regVec_0 = regVec_3746;
      end
      12'b111010100011 : begin
        _zz__zz_regVec_0 = regVec_3747;
      end
      12'b111010100100 : begin
        _zz__zz_regVec_0 = regVec_3748;
      end
      12'b111010100101 : begin
        _zz__zz_regVec_0 = regVec_3749;
      end
      12'b111010100110 : begin
        _zz__zz_regVec_0 = regVec_3750;
      end
      12'b111010100111 : begin
        _zz__zz_regVec_0 = regVec_3751;
      end
      12'b111010101000 : begin
        _zz__zz_regVec_0 = regVec_3752;
      end
      12'b111010101001 : begin
        _zz__zz_regVec_0 = regVec_3753;
      end
      12'b111010101010 : begin
        _zz__zz_regVec_0 = regVec_3754;
      end
      12'b111010101011 : begin
        _zz__zz_regVec_0 = regVec_3755;
      end
      12'b111010101100 : begin
        _zz__zz_regVec_0 = regVec_3756;
      end
      12'b111010101101 : begin
        _zz__zz_regVec_0 = regVec_3757;
      end
      12'b111010101110 : begin
        _zz__zz_regVec_0 = regVec_3758;
      end
      12'b111010101111 : begin
        _zz__zz_regVec_0 = regVec_3759;
      end
      12'b111010110000 : begin
        _zz__zz_regVec_0 = regVec_3760;
      end
      12'b111010110001 : begin
        _zz__zz_regVec_0 = regVec_3761;
      end
      12'b111010110010 : begin
        _zz__zz_regVec_0 = regVec_3762;
      end
      12'b111010110011 : begin
        _zz__zz_regVec_0 = regVec_3763;
      end
      12'b111010110100 : begin
        _zz__zz_regVec_0 = regVec_3764;
      end
      12'b111010110101 : begin
        _zz__zz_regVec_0 = regVec_3765;
      end
      12'b111010110110 : begin
        _zz__zz_regVec_0 = regVec_3766;
      end
      12'b111010110111 : begin
        _zz__zz_regVec_0 = regVec_3767;
      end
      12'b111010111000 : begin
        _zz__zz_regVec_0 = regVec_3768;
      end
      12'b111010111001 : begin
        _zz__zz_regVec_0 = regVec_3769;
      end
      12'b111010111010 : begin
        _zz__zz_regVec_0 = regVec_3770;
      end
      12'b111010111011 : begin
        _zz__zz_regVec_0 = regVec_3771;
      end
      12'b111010111100 : begin
        _zz__zz_regVec_0 = regVec_3772;
      end
      12'b111010111101 : begin
        _zz__zz_regVec_0 = regVec_3773;
      end
      12'b111010111110 : begin
        _zz__zz_regVec_0 = regVec_3774;
      end
      12'b111010111111 : begin
        _zz__zz_regVec_0 = regVec_3775;
      end
      12'b111011000000 : begin
        _zz__zz_regVec_0 = regVec_3776;
      end
      12'b111011000001 : begin
        _zz__zz_regVec_0 = regVec_3777;
      end
      12'b111011000010 : begin
        _zz__zz_regVec_0 = regVec_3778;
      end
      12'b111011000011 : begin
        _zz__zz_regVec_0 = regVec_3779;
      end
      12'b111011000100 : begin
        _zz__zz_regVec_0 = regVec_3780;
      end
      12'b111011000101 : begin
        _zz__zz_regVec_0 = regVec_3781;
      end
      12'b111011000110 : begin
        _zz__zz_regVec_0 = regVec_3782;
      end
      12'b111011000111 : begin
        _zz__zz_regVec_0 = regVec_3783;
      end
      12'b111011001000 : begin
        _zz__zz_regVec_0 = regVec_3784;
      end
      12'b111011001001 : begin
        _zz__zz_regVec_0 = regVec_3785;
      end
      12'b111011001010 : begin
        _zz__zz_regVec_0 = regVec_3786;
      end
      12'b111011001011 : begin
        _zz__zz_regVec_0 = regVec_3787;
      end
      12'b111011001100 : begin
        _zz__zz_regVec_0 = regVec_3788;
      end
      12'b111011001101 : begin
        _zz__zz_regVec_0 = regVec_3789;
      end
      12'b111011001110 : begin
        _zz__zz_regVec_0 = regVec_3790;
      end
      12'b111011001111 : begin
        _zz__zz_regVec_0 = regVec_3791;
      end
      12'b111011010000 : begin
        _zz__zz_regVec_0 = regVec_3792;
      end
      12'b111011010001 : begin
        _zz__zz_regVec_0 = regVec_3793;
      end
      12'b111011010010 : begin
        _zz__zz_regVec_0 = regVec_3794;
      end
      12'b111011010011 : begin
        _zz__zz_regVec_0 = regVec_3795;
      end
      12'b111011010100 : begin
        _zz__zz_regVec_0 = regVec_3796;
      end
      12'b111011010101 : begin
        _zz__zz_regVec_0 = regVec_3797;
      end
      12'b111011010110 : begin
        _zz__zz_regVec_0 = regVec_3798;
      end
      12'b111011010111 : begin
        _zz__zz_regVec_0 = regVec_3799;
      end
      12'b111011011000 : begin
        _zz__zz_regVec_0 = regVec_3800;
      end
      12'b111011011001 : begin
        _zz__zz_regVec_0 = regVec_3801;
      end
      12'b111011011010 : begin
        _zz__zz_regVec_0 = regVec_3802;
      end
      12'b111011011011 : begin
        _zz__zz_regVec_0 = regVec_3803;
      end
      12'b111011011100 : begin
        _zz__zz_regVec_0 = regVec_3804;
      end
      12'b111011011101 : begin
        _zz__zz_regVec_0 = regVec_3805;
      end
      12'b111011011110 : begin
        _zz__zz_regVec_0 = regVec_3806;
      end
      12'b111011011111 : begin
        _zz__zz_regVec_0 = regVec_3807;
      end
      12'b111011100000 : begin
        _zz__zz_regVec_0 = regVec_3808;
      end
      12'b111011100001 : begin
        _zz__zz_regVec_0 = regVec_3809;
      end
      12'b111011100010 : begin
        _zz__zz_regVec_0 = regVec_3810;
      end
      12'b111011100011 : begin
        _zz__zz_regVec_0 = regVec_3811;
      end
      12'b111011100100 : begin
        _zz__zz_regVec_0 = regVec_3812;
      end
      12'b111011100101 : begin
        _zz__zz_regVec_0 = regVec_3813;
      end
      12'b111011100110 : begin
        _zz__zz_regVec_0 = regVec_3814;
      end
      12'b111011100111 : begin
        _zz__zz_regVec_0 = regVec_3815;
      end
      12'b111011101000 : begin
        _zz__zz_regVec_0 = regVec_3816;
      end
      12'b111011101001 : begin
        _zz__zz_regVec_0 = regVec_3817;
      end
      12'b111011101010 : begin
        _zz__zz_regVec_0 = regVec_3818;
      end
      12'b111011101011 : begin
        _zz__zz_regVec_0 = regVec_3819;
      end
      12'b111011101100 : begin
        _zz__zz_regVec_0 = regVec_3820;
      end
      12'b111011101101 : begin
        _zz__zz_regVec_0 = regVec_3821;
      end
      12'b111011101110 : begin
        _zz__zz_regVec_0 = regVec_3822;
      end
      12'b111011101111 : begin
        _zz__zz_regVec_0 = regVec_3823;
      end
      12'b111011110000 : begin
        _zz__zz_regVec_0 = regVec_3824;
      end
      12'b111011110001 : begin
        _zz__zz_regVec_0 = regVec_3825;
      end
      12'b111011110010 : begin
        _zz__zz_regVec_0 = regVec_3826;
      end
      12'b111011110011 : begin
        _zz__zz_regVec_0 = regVec_3827;
      end
      12'b111011110100 : begin
        _zz__zz_regVec_0 = regVec_3828;
      end
      12'b111011110101 : begin
        _zz__zz_regVec_0 = regVec_3829;
      end
      12'b111011110110 : begin
        _zz__zz_regVec_0 = regVec_3830;
      end
      12'b111011110111 : begin
        _zz__zz_regVec_0 = regVec_3831;
      end
      12'b111011111000 : begin
        _zz__zz_regVec_0 = regVec_3832;
      end
      12'b111011111001 : begin
        _zz__zz_regVec_0 = regVec_3833;
      end
      12'b111011111010 : begin
        _zz__zz_regVec_0 = regVec_3834;
      end
      12'b111011111011 : begin
        _zz__zz_regVec_0 = regVec_3835;
      end
      12'b111011111100 : begin
        _zz__zz_regVec_0 = regVec_3836;
      end
      12'b111011111101 : begin
        _zz__zz_regVec_0 = regVec_3837;
      end
      12'b111011111110 : begin
        _zz__zz_regVec_0 = regVec_3838;
      end
      12'b111011111111 : begin
        _zz__zz_regVec_0 = regVec_3839;
      end
      12'b111100000000 : begin
        _zz__zz_regVec_0 = regVec_3840;
      end
      12'b111100000001 : begin
        _zz__zz_regVec_0 = regVec_3841;
      end
      12'b111100000010 : begin
        _zz__zz_regVec_0 = regVec_3842;
      end
      12'b111100000011 : begin
        _zz__zz_regVec_0 = regVec_3843;
      end
      12'b111100000100 : begin
        _zz__zz_regVec_0 = regVec_3844;
      end
      12'b111100000101 : begin
        _zz__zz_regVec_0 = regVec_3845;
      end
      12'b111100000110 : begin
        _zz__zz_regVec_0 = regVec_3846;
      end
      12'b111100000111 : begin
        _zz__zz_regVec_0 = regVec_3847;
      end
      12'b111100001000 : begin
        _zz__zz_regVec_0 = regVec_3848;
      end
      12'b111100001001 : begin
        _zz__zz_regVec_0 = regVec_3849;
      end
      12'b111100001010 : begin
        _zz__zz_regVec_0 = regVec_3850;
      end
      12'b111100001011 : begin
        _zz__zz_regVec_0 = regVec_3851;
      end
      12'b111100001100 : begin
        _zz__zz_regVec_0 = regVec_3852;
      end
      12'b111100001101 : begin
        _zz__zz_regVec_0 = regVec_3853;
      end
      12'b111100001110 : begin
        _zz__zz_regVec_0 = regVec_3854;
      end
      12'b111100001111 : begin
        _zz__zz_regVec_0 = regVec_3855;
      end
      12'b111100010000 : begin
        _zz__zz_regVec_0 = regVec_3856;
      end
      12'b111100010001 : begin
        _zz__zz_regVec_0 = regVec_3857;
      end
      12'b111100010010 : begin
        _zz__zz_regVec_0 = regVec_3858;
      end
      12'b111100010011 : begin
        _zz__zz_regVec_0 = regVec_3859;
      end
      12'b111100010100 : begin
        _zz__zz_regVec_0 = regVec_3860;
      end
      12'b111100010101 : begin
        _zz__zz_regVec_0 = regVec_3861;
      end
      12'b111100010110 : begin
        _zz__zz_regVec_0 = regVec_3862;
      end
      12'b111100010111 : begin
        _zz__zz_regVec_0 = regVec_3863;
      end
      12'b111100011000 : begin
        _zz__zz_regVec_0 = regVec_3864;
      end
      12'b111100011001 : begin
        _zz__zz_regVec_0 = regVec_3865;
      end
      12'b111100011010 : begin
        _zz__zz_regVec_0 = regVec_3866;
      end
      12'b111100011011 : begin
        _zz__zz_regVec_0 = regVec_3867;
      end
      12'b111100011100 : begin
        _zz__zz_regVec_0 = regVec_3868;
      end
      12'b111100011101 : begin
        _zz__zz_regVec_0 = regVec_3869;
      end
      12'b111100011110 : begin
        _zz__zz_regVec_0 = regVec_3870;
      end
      12'b111100011111 : begin
        _zz__zz_regVec_0 = regVec_3871;
      end
      12'b111100100000 : begin
        _zz__zz_regVec_0 = regVec_3872;
      end
      12'b111100100001 : begin
        _zz__zz_regVec_0 = regVec_3873;
      end
      12'b111100100010 : begin
        _zz__zz_regVec_0 = regVec_3874;
      end
      12'b111100100011 : begin
        _zz__zz_regVec_0 = regVec_3875;
      end
      12'b111100100100 : begin
        _zz__zz_regVec_0 = regVec_3876;
      end
      12'b111100100101 : begin
        _zz__zz_regVec_0 = regVec_3877;
      end
      12'b111100100110 : begin
        _zz__zz_regVec_0 = regVec_3878;
      end
      12'b111100100111 : begin
        _zz__zz_regVec_0 = regVec_3879;
      end
      12'b111100101000 : begin
        _zz__zz_regVec_0 = regVec_3880;
      end
      12'b111100101001 : begin
        _zz__zz_regVec_0 = regVec_3881;
      end
      12'b111100101010 : begin
        _zz__zz_regVec_0 = regVec_3882;
      end
      12'b111100101011 : begin
        _zz__zz_regVec_0 = regVec_3883;
      end
      12'b111100101100 : begin
        _zz__zz_regVec_0 = regVec_3884;
      end
      12'b111100101101 : begin
        _zz__zz_regVec_0 = regVec_3885;
      end
      12'b111100101110 : begin
        _zz__zz_regVec_0 = regVec_3886;
      end
      12'b111100101111 : begin
        _zz__zz_regVec_0 = regVec_3887;
      end
      12'b111100110000 : begin
        _zz__zz_regVec_0 = regVec_3888;
      end
      12'b111100110001 : begin
        _zz__zz_regVec_0 = regVec_3889;
      end
      12'b111100110010 : begin
        _zz__zz_regVec_0 = regVec_3890;
      end
      12'b111100110011 : begin
        _zz__zz_regVec_0 = regVec_3891;
      end
      12'b111100110100 : begin
        _zz__zz_regVec_0 = regVec_3892;
      end
      12'b111100110101 : begin
        _zz__zz_regVec_0 = regVec_3893;
      end
      12'b111100110110 : begin
        _zz__zz_regVec_0 = regVec_3894;
      end
      12'b111100110111 : begin
        _zz__zz_regVec_0 = regVec_3895;
      end
      12'b111100111000 : begin
        _zz__zz_regVec_0 = regVec_3896;
      end
      12'b111100111001 : begin
        _zz__zz_regVec_0 = regVec_3897;
      end
      12'b111100111010 : begin
        _zz__zz_regVec_0 = regVec_3898;
      end
      12'b111100111011 : begin
        _zz__zz_regVec_0 = regVec_3899;
      end
      12'b111100111100 : begin
        _zz__zz_regVec_0 = regVec_3900;
      end
      12'b111100111101 : begin
        _zz__zz_regVec_0 = regVec_3901;
      end
      12'b111100111110 : begin
        _zz__zz_regVec_0 = regVec_3902;
      end
      12'b111100111111 : begin
        _zz__zz_regVec_0 = regVec_3903;
      end
      12'b111101000000 : begin
        _zz__zz_regVec_0 = regVec_3904;
      end
      12'b111101000001 : begin
        _zz__zz_regVec_0 = regVec_3905;
      end
      12'b111101000010 : begin
        _zz__zz_regVec_0 = regVec_3906;
      end
      12'b111101000011 : begin
        _zz__zz_regVec_0 = regVec_3907;
      end
      12'b111101000100 : begin
        _zz__zz_regVec_0 = regVec_3908;
      end
      12'b111101000101 : begin
        _zz__zz_regVec_0 = regVec_3909;
      end
      12'b111101000110 : begin
        _zz__zz_regVec_0 = regVec_3910;
      end
      12'b111101000111 : begin
        _zz__zz_regVec_0 = regVec_3911;
      end
      12'b111101001000 : begin
        _zz__zz_regVec_0 = regVec_3912;
      end
      12'b111101001001 : begin
        _zz__zz_regVec_0 = regVec_3913;
      end
      12'b111101001010 : begin
        _zz__zz_regVec_0 = regVec_3914;
      end
      12'b111101001011 : begin
        _zz__zz_regVec_0 = regVec_3915;
      end
      12'b111101001100 : begin
        _zz__zz_regVec_0 = regVec_3916;
      end
      12'b111101001101 : begin
        _zz__zz_regVec_0 = regVec_3917;
      end
      12'b111101001110 : begin
        _zz__zz_regVec_0 = regVec_3918;
      end
      12'b111101001111 : begin
        _zz__zz_regVec_0 = regVec_3919;
      end
      12'b111101010000 : begin
        _zz__zz_regVec_0 = regVec_3920;
      end
      12'b111101010001 : begin
        _zz__zz_regVec_0 = regVec_3921;
      end
      12'b111101010010 : begin
        _zz__zz_regVec_0 = regVec_3922;
      end
      12'b111101010011 : begin
        _zz__zz_regVec_0 = regVec_3923;
      end
      12'b111101010100 : begin
        _zz__zz_regVec_0 = regVec_3924;
      end
      12'b111101010101 : begin
        _zz__zz_regVec_0 = regVec_3925;
      end
      12'b111101010110 : begin
        _zz__zz_regVec_0 = regVec_3926;
      end
      12'b111101010111 : begin
        _zz__zz_regVec_0 = regVec_3927;
      end
      12'b111101011000 : begin
        _zz__zz_regVec_0 = regVec_3928;
      end
      12'b111101011001 : begin
        _zz__zz_regVec_0 = regVec_3929;
      end
      12'b111101011010 : begin
        _zz__zz_regVec_0 = regVec_3930;
      end
      12'b111101011011 : begin
        _zz__zz_regVec_0 = regVec_3931;
      end
      12'b111101011100 : begin
        _zz__zz_regVec_0 = regVec_3932;
      end
      12'b111101011101 : begin
        _zz__zz_regVec_0 = regVec_3933;
      end
      12'b111101011110 : begin
        _zz__zz_regVec_0 = regVec_3934;
      end
      12'b111101011111 : begin
        _zz__zz_regVec_0 = regVec_3935;
      end
      12'b111101100000 : begin
        _zz__zz_regVec_0 = regVec_3936;
      end
      12'b111101100001 : begin
        _zz__zz_regVec_0 = regVec_3937;
      end
      12'b111101100010 : begin
        _zz__zz_regVec_0 = regVec_3938;
      end
      12'b111101100011 : begin
        _zz__zz_regVec_0 = regVec_3939;
      end
      12'b111101100100 : begin
        _zz__zz_regVec_0 = regVec_3940;
      end
      12'b111101100101 : begin
        _zz__zz_regVec_0 = regVec_3941;
      end
      12'b111101100110 : begin
        _zz__zz_regVec_0 = regVec_3942;
      end
      12'b111101100111 : begin
        _zz__zz_regVec_0 = regVec_3943;
      end
      12'b111101101000 : begin
        _zz__zz_regVec_0 = regVec_3944;
      end
      12'b111101101001 : begin
        _zz__zz_regVec_0 = regVec_3945;
      end
      12'b111101101010 : begin
        _zz__zz_regVec_0 = regVec_3946;
      end
      12'b111101101011 : begin
        _zz__zz_regVec_0 = regVec_3947;
      end
      12'b111101101100 : begin
        _zz__zz_regVec_0 = regVec_3948;
      end
      12'b111101101101 : begin
        _zz__zz_regVec_0 = regVec_3949;
      end
      12'b111101101110 : begin
        _zz__zz_regVec_0 = regVec_3950;
      end
      12'b111101101111 : begin
        _zz__zz_regVec_0 = regVec_3951;
      end
      12'b111101110000 : begin
        _zz__zz_regVec_0 = regVec_3952;
      end
      12'b111101110001 : begin
        _zz__zz_regVec_0 = regVec_3953;
      end
      12'b111101110010 : begin
        _zz__zz_regVec_0 = regVec_3954;
      end
      12'b111101110011 : begin
        _zz__zz_regVec_0 = regVec_3955;
      end
      12'b111101110100 : begin
        _zz__zz_regVec_0 = regVec_3956;
      end
      12'b111101110101 : begin
        _zz__zz_regVec_0 = regVec_3957;
      end
      12'b111101110110 : begin
        _zz__zz_regVec_0 = regVec_3958;
      end
      12'b111101110111 : begin
        _zz__zz_regVec_0 = regVec_3959;
      end
      12'b111101111000 : begin
        _zz__zz_regVec_0 = regVec_3960;
      end
      12'b111101111001 : begin
        _zz__zz_regVec_0 = regVec_3961;
      end
      12'b111101111010 : begin
        _zz__zz_regVec_0 = regVec_3962;
      end
      12'b111101111011 : begin
        _zz__zz_regVec_0 = regVec_3963;
      end
      12'b111101111100 : begin
        _zz__zz_regVec_0 = regVec_3964;
      end
      12'b111101111101 : begin
        _zz__zz_regVec_0 = regVec_3965;
      end
      12'b111101111110 : begin
        _zz__zz_regVec_0 = regVec_3966;
      end
      12'b111101111111 : begin
        _zz__zz_regVec_0 = regVec_3967;
      end
      12'b111110000000 : begin
        _zz__zz_regVec_0 = regVec_3968;
      end
      12'b111110000001 : begin
        _zz__zz_regVec_0 = regVec_3969;
      end
      12'b111110000010 : begin
        _zz__zz_regVec_0 = regVec_3970;
      end
      12'b111110000011 : begin
        _zz__zz_regVec_0 = regVec_3971;
      end
      12'b111110000100 : begin
        _zz__zz_regVec_0 = regVec_3972;
      end
      12'b111110000101 : begin
        _zz__zz_regVec_0 = regVec_3973;
      end
      12'b111110000110 : begin
        _zz__zz_regVec_0 = regVec_3974;
      end
      12'b111110000111 : begin
        _zz__zz_regVec_0 = regVec_3975;
      end
      12'b111110001000 : begin
        _zz__zz_regVec_0 = regVec_3976;
      end
      12'b111110001001 : begin
        _zz__zz_regVec_0 = regVec_3977;
      end
      12'b111110001010 : begin
        _zz__zz_regVec_0 = regVec_3978;
      end
      12'b111110001011 : begin
        _zz__zz_regVec_0 = regVec_3979;
      end
      12'b111110001100 : begin
        _zz__zz_regVec_0 = regVec_3980;
      end
      12'b111110001101 : begin
        _zz__zz_regVec_0 = regVec_3981;
      end
      12'b111110001110 : begin
        _zz__zz_regVec_0 = regVec_3982;
      end
      12'b111110001111 : begin
        _zz__zz_regVec_0 = regVec_3983;
      end
      12'b111110010000 : begin
        _zz__zz_regVec_0 = regVec_3984;
      end
      12'b111110010001 : begin
        _zz__zz_regVec_0 = regVec_3985;
      end
      12'b111110010010 : begin
        _zz__zz_regVec_0 = regVec_3986;
      end
      12'b111110010011 : begin
        _zz__zz_regVec_0 = regVec_3987;
      end
      12'b111110010100 : begin
        _zz__zz_regVec_0 = regVec_3988;
      end
      12'b111110010101 : begin
        _zz__zz_regVec_0 = regVec_3989;
      end
      12'b111110010110 : begin
        _zz__zz_regVec_0 = regVec_3990;
      end
      12'b111110010111 : begin
        _zz__zz_regVec_0 = regVec_3991;
      end
      12'b111110011000 : begin
        _zz__zz_regVec_0 = regVec_3992;
      end
      12'b111110011001 : begin
        _zz__zz_regVec_0 = regVec_3993;
      end
      12'b111110011010 : begin
        _zz__zz_regVec_0 = regVec_3994;
      end
      12'b111110011011 : begin
        _zz__zz_regVec_0 = regVec_3995;
      end
      12'b111110011100 : begin
        _zz__zz_regVec_0 = regVec_3996;
      end
      12'b111110011101 : begin
        _zz__zz_regVec_0 = regVec_3997;
      end
      12'b111110011110 : begin
        _zz__zz_regVec_0 = regVec_3998;
      end
      12'b111110011111 : begin
        _zz__zz_regVec_0 = regVec_3999;
      end
      12'b111110100000 : begin
        _zz__zz_regVec_0 = regVec_4000;
      end
      12'b111110100001 : begin
        _zz__zz_regVec_0 = regVec_4001;
      end
      12'b111110100010 : begin
        _zz__zz_regVec_0 = regVec_4002;
      end
      12'b111110100011 : begin
        _zz__zz_regVec_0 = regVec_4003;
      end
      12'b111110100100 : begin
        _zz__zz_regVec_0 = regVec_4004;
      end
      12'b111110100101 : begin
        _zz__zz_regVec_0 = regVec_4005;
      end
      12'b111110100110 : begin
        _zz__zz_regVec_0 = regVec_4006;
      end
      12'b111110100111 : begin
        _zz__zz_regVec_0 = regVec_4007;
      end
      12'b111110101000 : begin
        _zz__zz_regVec_0 = regVec_4008;
      end
      12'b111110101001 : begin
        _zz__zz_regVec_0 = regVec_4009;
      end
      12'b111110101010 : begin
        _zz__zz_regVec_0 = regVec_4010;
      end
      12'b111110101011 : begin
        _zz__zz_regVec_0 = regVec_4011;
      end
      12'b111110101100 : begin
        _zz__zz_regVec_0 = regVec_4012;
      end
      12'b111110101101 : begin
        _zz__zz_regVec_0 = regVec_4013;
      end
      12'b111110101110 : begin
        _zz__zz_regVec_0 = regVec_4014;
      end
      12'b111110101111 : begin
        _zz__zz_regVec_0 = regVec_4015;
      end
      12'b111110110000 : begin
        _zz__zz_regVec_0 = regVec_4016;
      end
      12'b111110110001 : begin
        _zz__zz_regVec_0 = regVec_4017;
      end
      12'b111110110010 : begin
        _zz__zz_regVec_0 = regVec_4018;
      end
      12'b111110110011 : begin
        _zz__zz_regVec_0 = regVec_4019;
      end
      12'b111110110100 : begin
        _zz__zz_regVec_0 = regVec_4020;
      end
      12'b111110110101 : begin
        _zz__zz_regVec_0 = regVec_4021;
      end
      12'b111110110110 : begin
        _zz__zz_regVec_0 = regVec_4022;
      end
      12'b111110110111 : begin
        _zz__zz_regVec_0 = regVec_4023;
      end
      12'b111110111000 : begin
        _zz__zz_regVec_0 = regVec_4024;
      end
      12'b111110111001 : begin
        _zz__zz_regVec_0 = regVec_4025;
      end
      12'b111110111010 : begin
        _zz__zz_regVec_0 = regVec_4026;
      end
      12'b111110111011 : begin
        _zz__zz_regVec_0 = regVec_4027;
      end
      12'b111110111100 : begin
        _zz__zz_regVec_0 = regVec_4028;
      end
      12'b111110111101 : begin
        _zz__zz_regVec_0 = regVec_4029;
      end
      12'b111110111110 : begin
        _zz__zz_regVec_0 = regVec_4030;
      end
      12'b111110111111 : begin
        _zz__zz_regVec_0 = regVec_4031;
      end
      12'b111111000000 : begin
        _zz__zz_regVec_0 = regVec_4032;
      end
      12'b111111000001 : begin
        _zz__zz_regVec_0 = regVec_4033;
      end
      12'b111111000010 : begin
        _zz__zz_regVec_0 = regVec_4034;
      end
      12'b111111000011 : begin
        _zz__zz_regVec_0 = regVec_4035;
      end
      12'b111111000100 : begin
        _zz__zz_regVec_0 = regVec_4036;
      end
      12'b111111000101 : begin
        _zz__zz_regVec_0 = regVec_4037;
      end
      12'b111111000110 : begin
        _zz__zz_regVec_0 = regVec_4038;
      end
      12'b111111000111 : begin
        _zz__zz_regVec_0 = regVec_4039;
      end
      12'b111111001000 : begin
        _zz__zz_regVec_0 = regVec_4040;
      end
      12'b111111001001 : begin
        _zz__zz_regVec_0 = regVec_4041;
      end
      12'b111111001010 : begin
        _zz__zz_regVec_0 = regVec_4042;
      end
      12'b111111001011 : begin
        _zz__zz_regVec_0 = regVec_4043;
      end
      12'b111111001100 : begin
        _zz__zz_regVec_0 = regVec_4044;
      end
      12'b111111001101 : begin
        _zz__zz_regVec_0 = regVec_4045;
      end
      12'b111111001110 : begin
        _zz__zz_regVec_0 = regVec_4046;
      end
      12'b111111001111 : begin
        _zz__zz_regVec_0 = regVec_4047;
      end
      12'b111111010000 : begin
        _zz__zz_regVec_0 = regVec_4048;
      end
      12'b111111010001 : begin
        _zz__zz_regVec_0 = regVec_4049;
      end
      12'b111111010010 : begin
        _zz__zz_regVec_0 = regVec_4050;
      end
      12'b111111010011 : begin
        _zz__zz_regVec_0 = regVec_4051;
      end
      12'b111111010100 : begin
        _zz__zz_regVec_0 = regVec_4052;
      end
      12'b111111010101 : begin
        _zz__zz_regVec_0 = regVec_4053;
      end
      12'b111111010110 : begin
        _zz__zz_regVec_0 = regVec_4054;
      end
      12'b111111010111 : begin
        _zz__zz_regVec_0 = regVec_4055;
      end
      12'b111111011000 : begin
        _zz__zz_regVec_0 = regVec_4056;
      end
      12'b111111011001 : begin
        _zz__zz_regVec_0 = regVec_4057;
      end
      12'b111111011010 : begin
        _zz__zz_regVec_0 = regVec_4058;
      end
      12'b111111011011 : begin
        _zz__zz_regVec_0 = regVec_4059;
      end
      12'b111111011100 : begin
        _zz__zz_regVec_0 = regVec_4060;
      end
      12'b111111011101 : begin
        _zz__zz_regVec_0 = regVec_4061;
      end
      12'b111111011110 : begin
        _zz__zz_regVec_0 = regVec_4062;
      end
      12'b111111011111 : begin
        _zz__zz_regVec_0 = regVec_4063;
      end
      12'b111111100000 : begin
        _zz__zz_regVec_0 = regVec_4064;
      end
      12'b111111100001 : begin
        _zz__zz_regVec_0 = regVec_4065;
      end
      12'b111111100010 : begin
        _zz__zz_regVec_0 = regVec_4066;
      end
      12'b111111100011 : begin
        _zz__zz_regVec_0 = regVec_4067;
      end
      12'b111111100100 : begin
        _zz__zz_regVec_0 = regVec_4068;
      end
      12'b111111100101 : begin
        _zz__zz_regVec_0 = regVec_4069;
      end
      12'b111111100110 : begin
        _zz__zz_regVec_0 = regVec_4070;
      end
      12'b111111100111 : begin
        _zz__zz_regVec_0 = regVec_4071;
      end
      12'b111111101000 : begin
        _zz__zz_regVec_0 = regVec_4072;
      end
      12'b111111101001 : begin
        _zz__zz_regVec_0 = regVec_4073;
      end
      12'b111111101010 : begin
        _zz__zz_regVec_0 = regVec_4074;
      end
      12'b111111101011 : begin
        _zz__zz_regVec_0 = regVec_4075;
      end
      12'b111111101100 : begin
        _zz__zz_regVec_0 = regVec_4076;
      end
      12'b111111101101 : begin
        _zz__zz_regVec_0 = regVec_4077;
      end
      12'b111111101110 : begin
        _zz__zz_regVec_0 = regVec_4078;
      end
      12'b111111101111 : begin
        _zz__zz_regVec_0 = regVec_4079;
      end
      12'b111111110000 : begin
        _zz__zz_regVec_0 = regVec_4080;
      end
      12'b111111110001 : begin
        _zz__zz_regVec_0 = regVec_4081;
      end
      12'b111111110010 : begin
        _zz__zz_regVec_0 = regVec_4082;
      end
      12'b111111110011 : begin
        _zz__zz_regVec_0 = regVec_4083;
      end
      12'b111111110100 : begin
        _zz__zz_regVec_0 = regVec_4084;
      end
      12'b111111110101 : begin
        _zz__zz_regVec_0 = regVec_4085;
      end
      12'b111111110110 : begin
        _zz__zz_regVec_0 = regVec_4086;
      end
      12'b111111110111 : begin
        _zz__zz_regVec_0 = regVec_4087;
      end
      12'b111111111000 : begin
        _zz__zz_regVec_0 = regVec_4088;
      end
      12'b111111111001 : begin
        _zz__zz_regVec_0 = regVec_4089;
      end
      12'b111111111010 : begin
        _zz__zz_regVec_0 = regVec_4090;
      end
      12'b111111111011 : begin
        _zz__zz_regVec_0 = regVec_4091;
      end
      12'b111111111100 : begin
        _zz__zz_regVec_0 = regVec_4092;
      end
      12'b111111111101 : begin
        _zz__zz_regVec_0 = regVec_4093;
      end
      12'b111111111110 : begin
        _zz__zz_regVec_0 = regVec_4094;
      end
      default : begin
        _zz__zz_regVec_0 = regVec_4095;
      end
    endcase
  end

  always @(*) begin
    case(regAwAddr)
      12'b000000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_0;
      end
      12'b000000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1;
      end
      12'b000000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2;
      end
      12'b000000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3;
      end
      12'b000000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4;
      end
      12'b000000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_5;
      end
      12'b000000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_6;
      end
      12'b000000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_7;
      end
      12'b000000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_8;
      end
      12'b000000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_9;
      end
      12'b000000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_10;
      end
      12'b000000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_11;
      end
      12'b000000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_12;
      end
      12'b000000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_13;
      end
      12'b000000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_14;
      end
      12'b000000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_15;
      end
      12'b000000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_16;
      end
      12'b000000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_17;
      end
      12'b000000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_18;
      end
      12'b000000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_19;
      end
      12'b000000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_20;
      end
      12'b000000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_21;
      end
      12'b000000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_22;
      end
      12'b000000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_23;
      end
      12'b000000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_24;
      end
      12'b000000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_25;
      end
      12'b000000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_26;
      end
      12'b000000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_27;
      end
      12'b000000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_28;
      end
      12'b000000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_29;
      end
      12'b000000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_30;
      end
      12'b000000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_31;
      end
      12'b000000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_32;
      end
      12'b000000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_33;
      end
      12'b000000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_34;
      end
      12'b000000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_35;
      end
      12'b000000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_36;
      end
      12'b000000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_37;
      end
      12'b000000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_38;
      end
      12'b000000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_39;
      end
      12'b000000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_40;
      end
      12'b000000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_41;
      end
      12'b000000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_42;
      end
      12'b000000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_43;
      end
      12'b000000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_44;
      end
      12'b000000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_45;
      end
      12'b000000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_46;
      end
      12'b000000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_47;
      end
      12'b000000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_48;
      end
      12'b000000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_49;
      end
      12'b000000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_50;
      end
      12'b000000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_51;
      end
      12'b000000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_52;
      end
      12'b000000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_53;
      end
      12'b000000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_54;
      end
      12'b000000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_55;
      end
      12'b000000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_56;
      end
      12'b000000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_57;
      end
      12'b000000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_58;
      end
      12'b000000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_59;
      end
      12'b000000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_60;
      end
      12'b000000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_61;
      end
      12'b000000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_62;
      end
      12'b000000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_63;
      end
      12'b000001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_64;
      end
      12'b000001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_65;
      end
      12'b000001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_66;
      end
      12'b000001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_67;
      end
      12'b000001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_68;
      end
      12'b000001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_69;
      end
      12'b000001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_70;
      end
      12'b000001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_71;
      end
      12'b000001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_72;
      end
      12'b000001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_73;
      end
      12'b000001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_74;
      end
      12'b000001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_75;
      end
      12'b000001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_76;
      end
      12'b000001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_77;
      end
      12'b000001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_78;
      end
      12'b000001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_79;
      end
      12'b000001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_80;
      end
      12'b000001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_81;
      end
      12'b000001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_82;
      end
      12'b000001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_83;
      end
      12'b000001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_84;
      end
      12'b000001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_85;
      end
      12'b000001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_86;
      end
      12'b000001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_87;
      end
      12'b000001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_88;
      end
      12'b000001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_89;
      end
      12'b000001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_90;
      end
      12'b000001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_91;
      end
      12'b000001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_92;
      end
      12'b000001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_93;
      end
      12'b000001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_94;
      end
      12'b000001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_95;
      end
      12'b000001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_96;
      end
      12'b000001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_97;
      end
      12'b000001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_98;
      end
      12'b000001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_99;
      end
      12'b000001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_100;
      end
      12'b000001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_101;
      end
      12'b000001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_102;
      end
      12'b000001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_103;
      end
      12'b000001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_104;
      end
      12'b000001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_105;
      end
      12'b000001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_106;
      end
      12'b000001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_107;
      end
      12'b000001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_108;
      end
      12'b000001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_109;
      end
      12'b000001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_110;
      end
      12'b000001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_111;
      end
      12'b000001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_112;
      end
      12'b000001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_113;
      end
      12'b000001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_114;
      end
      12'b000001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_115;
      end
      12'b000001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_116;
      end
      12'b000001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_117;
      end
      12'b000001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_118;
      end
      12'b000001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_119;
      end
      12'b000001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_120;
      end
      12'b000001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_121;
      end
      12'b000001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_122;
      end
      12'b000001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_123;
      end
      12'b000001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_124;
      end
      12'b000001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_125;
      end
      12'b000001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_126;
      end
      12'b000001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_127;
      end
      12'b000010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_128;
      end
      12'b000010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_129;
      end
      12'b000010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_130;
      end
      12'b000010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_131;
      end
      12'b000010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_132;
      end
      12'b000010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_133;
      end
      12'b000010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_134;
      end
      12'b000010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_135;
      end
      12'b000010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_136;
      end
      12'b000010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_137;
      end
      12'b000010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_138;
      end
      12'b000010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_139;
      end
      12'b000010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_140;
      end
      12'b000010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_141;
      end
      12'b000010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_142;
      end
      12'b000010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_143;
      end
      12'b000010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_144;
      end
      12'b000010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_145;
      end
      12'b000010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_146;
      end
      12'b000010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_147;
      end
      12'b000010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_148;
      end
      12'b000010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_149;
      end
      12'b000010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_150;
      end
      12'b000010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_151;
      end
      12'b000010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_152;
      end
      12'b000010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_153;
      end
      12'b000010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_154;
      end
      12'b000010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_155;
      end
      12'b000010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_156;
      end
      12'b000010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_157;
      end
      12'b000010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_158;
      end
      12'b000010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_159;
      end
      12'b000010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_160;
      end
      12'b000010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_161;
      end
      12'b000010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_162;
      end
      12'b000010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_163;
      end
      12'b000010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_164;
      end
      12'b000010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_165;
      end
      12'b000010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_166;
      end
      12'b000010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_167;
      end
      12'b000010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_168;
      end
      12'b000010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_169;
      end
      12'b000010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_170;
      end
      12'b000010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_171;
      end
      12'b000010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_172;
      end
      12'b000010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_173;
      end
      12'b000010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_174;
      end
      12'b000010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_175;
      end
      12'b000010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_176;
      end
      12'b000010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_177;
      end
      12'b000010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_178;
      end
      12'b000010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_179;
      end
      12'b000010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_180;
      end
      12'b000010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_181;
      end
      12'b000010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_182;
      end
      12'b000010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_183;
      end
      12'b000010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_184;
      end
      12'b000010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_185;
      end
      12'b000010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_186;
      end
      12'b000010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_187;
      end
      12'b000010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_188;
      end
      12'b000010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_189;
      end
      12'b000010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_190;
      end
      12'b000010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_191;
      end
      12'b000011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_192;
      end
      12'b000011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_193;
      end
      12'b000011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_194;
      end
      12'b000011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_195;
      end
      12'b000011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_196;
      end
      12'b000011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_197;
      end
      12'b000011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_198;
      end
      12'b000011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_199;
      end
      12'b000011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_200;
      end
      12'b000011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_201;
      end
      12'b000011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_202;
      end
      12'b000011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_203;
      end
      12'b000011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_204;
      end
      12'b000011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_205;
      end
      12'b000011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_206;
      end
      12'b000011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_207;
      end
      12'b000011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_208;
      end
      12'b000011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_209;
      end
      12'b000011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_210;
      end
      12'b000011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_211;
      end
      12'b000011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_212;
      end
      12'b000011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_213;
      end
      12'b000011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_214;
      end
      12'b000011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_215;
      end
      12'b000011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_216;
      end
      12'b000011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_217;
      end
      12'b000011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_218;
      end
      12'b000011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_219;
      end
      12'b000011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_220;
      end
      12'b000011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_221;
      end
      12'b000011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_222;
      end
      12'b000011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_223;
      end
      12'b000011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_224;
      end
      12'b000011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_225;
      end
      12'b000011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_226;
      end
      12'b000011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_227;
      end
      12'b000011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_228;
      end
      12'b000011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_229;
      end
      12'b000011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_230;
      end
      12'b000011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_231;
      end
      12'b000011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_232;
      end
      12'b000011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_233;
      end
      12'b000011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_234;
      end
      12'b000011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_235;
      end
      12'b000011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_236;
      end
      12'b000011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_237;
      end
      12'b000011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_238;
      end
      12'b000011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_239;
      end
      12'b000011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_240;
      end
      12'b000011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_241;
      end
      12'b000011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_242;
      end
      12'b000011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_243;
      end
      12'b000011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_244;
      end
      12'b000011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_245;
      end
      12'b000011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_246;
      end
      12'b000011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_247;
      end
      12'b000011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_248;
      end
      12'b000011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_249;
      end
      12'b000011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_250;
      end
      12'b000011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_251;
      end
      12'b000011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_252;
      end
      12'b000011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_253;
      end
      12'b000011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_254;
      end
      12'b000011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_255;
      end
      12'b000100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_256;
      end
      12'b000100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_257;
      end
      12'b000100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_258;
      end
      12'b000100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_259;
      end
      12'b000100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_260;
      end
      12'b000100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_261;
      end
      12'b000100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_262;
      end
      12'b000100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_263;
      end
      12'b000100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_264;
      end
      12'b000100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_265;
      end
      12'b000100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_266;
      end
      12'b000100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_267;
      end
      12'b000100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_268;
      end
      12'b000100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_269;
      end
      12'b000100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_270;
      end
      12'b000100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_271;
      end
      12'b000100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_272;
      end
      12'b000100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_273;
      end
      12'b000100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_274;
      end
      12'b000100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_275;
      end
      12'b000100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_276;
      end
      12'b000100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_277;
      end
      12'b000100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_278;
      end
      12'b000100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_279;
      end
      12'b000100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_280;
      end
      12'b000100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_281;
      end
      12'b000100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_282;
      end
      12'b000100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_283;
      end
      12'b000100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_284;
      end
      12'b000100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_285;
      end
      12'b000100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_286;
      end
      12'b000100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_287;
      end
      12'b000100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_288;
      end
      12'b000100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_289;
      end
      12'b000100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_290;
      end
      12'b000100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_291;
      end
      12'b000100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_292;
      end
      12'b000100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_293;
      end
      12'b000100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_294;
      end
      12'b000100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_295;
      end
      12'b000100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_296;
      end
      12'b000100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_297;
      end
      12'b000100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_298;
      end
      12'b000100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_299;
      end
      12'b000100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_300;
      end
      12'b000100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_301;
      end
      12'b000100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_302;
      end
      12'b000100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_303;
      end
      12'b000100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_304;
      end
      12'b000100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_305;
      end
      12'b000100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_306;
      end
      12'b000100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_307;
      end
      12'b000100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_308;
      end
      12'b000100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_309;
      end
      12'b000100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_310;
      end
      12'b000100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_311;
      end
      12'b000100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_312;
      end
      12'b000100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_313;
      end
      12'b000100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_314;
      end
      12'b000100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_315;
      end
      12'b000100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_316;
      end
      12'b000100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_317;
      end
      12'b000100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_318;
      end
      12'b000100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_319;
      end
      12'b000101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_320;
      end
      12'b000101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_321;
      end
      12'b000101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_322;
      end
      12'b000101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_323;
      end
      12'b000101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_324;
      end
      12'b000101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_325;
      end
      12'b000101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_326;
      end
      12'b000101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_327;
      end
      12'b000101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_328;
      end
      12'b000101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_329;
      end
      12'b000101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_330;
      end
      12'b000101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_331;
      end
      12'b000101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_332;
      end
      12'b000101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_333;
      end
      12'b000101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_334;
      end
      12'b000101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_335;
      end
      12'b000101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_336;
      end
      12'b000101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_337;
      end
      12'b000101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_338;
      end
      12'b000101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_339;
      end
      12'b000101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_340;
      end
      12'b000101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_341;
      end
      12'b000101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_342;
      end
      12'b000101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_343;
      end
      12'b000101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_344;
      end
      12'b000101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_345;
      end
      12'b000101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_346;
      end
      12'b000101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_347;
      end
      12'b000101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_348;
      end
      12'b000101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_349;
      end
      12'b000101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_350;
      end
      12'b000101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_351;
      end
      12'b000101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_352;
      end
      12'b000101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_353;
      end
      12'b000101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_354;
      end
      12'b000101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_355;
      end
      12'b000101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_356;
      end
      12'b000101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_357;
      end
      12'b000101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_358;
      end
      12'b000101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_359;
      end
      12'b000101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_360;
      end
      12'b000101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_361;
      end
      12'b000101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_362;
      end
      12'b000101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_363;
      end
      12'b000101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_364;
      end
      12'b000101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_365;
      end
      12'b000101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_366;
      end
      12'b000101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_367;
      end
      12'b000101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_368;
      end
      12'b000101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_369;
      end
      12'b000101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_370;
      end
      12'b000101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_371;
      end
      12'b000101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_372;
      end
      12'b000101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_373;
      end
      12'b000101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_374;
      end
      12'b000101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_375;
      end
      12'b000101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_376;
      end
      12'b000101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_377;
      end
      12'b000101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_378;
      end
      12'b000101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_379;
      end
      12'b000101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_380;
      end
      12'b000101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_381;
      end
      12'b000101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_382;
      end
      12'b000101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_383;
      end
      12'b000110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_384;
      end
      12'b000110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_385;
      end
      12'b000110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_386;
      end
      12'b000110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_387;
      end
      12'b000110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_388;
      end
      12'b000110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_389;
      end
      12'b000110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_390;
      end
      12'b000110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_391;
      end
      12'b000110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_392;
      end
      12'b000110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_393;
      end
      12'b000110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_394;
      end
      12'b000110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_395;
      end
      12'b000110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_396;
      end
      12'b000110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_397;
      end
      12'b000110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_398;
      end
      12'b000110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_399;
      end
      12'b000110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_400;
      end
      12'b000110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_401;
      end
      12'b000110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_402;
      end
      12'b000110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_403;
      end
      12'b000110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_404;
      end
      12'b000110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_405;
      end
      12'b000110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_406;
      end
      12'b000110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_407;
      end
      12'b000110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_408;
      end
      12'b000110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_409;
      end
      12'b000110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_410;
      end
      12'b000110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_411;
      end
      12'b000110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_412;
      end
      12'b000110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_413;
      end
      12'b000110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_414;
      end
      12'b000110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_415;
      end
      12'b000110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_416;
      end
      12'b000110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_417;
      end
      12'b000110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_418;
      end
      12'b000110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_419;
      end
      12'b000110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_420;
      end
      12'b000110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_421;
      end
      12'b000110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_422;
      end
      12'b000110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_423;
      end
      12'b000110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_424;
      end
      12'b000110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_425;
      end
      12'b000110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_426;
      end
      12'b000110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_427;
      end
      12'b000110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_428;
      end
      12'b000110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_429;
      end
      12'b000110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_430;
      end
      12'b000110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_431;
      end
      12'b000110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_432;
      end
      12'b000110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_433;
      end
      12'b000110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_434;
      end
      12'b000110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_435;
      end
      12'b000110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_436;
      end
      12'b000110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_437;
      end
      12'b000110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_438;
      end
      12'b000110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_439;
      end
      12'b000110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_440;
      end
      12'b000110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_441;
      end
      12'b000110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_442;
      end
      12'b000110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_443;
      end
      12'b000110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_444;
      end
      12'b000110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_445;
      end
      12'b000110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_446;
      end
      12'b000110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_447;
      end
      12'b000111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_448;
      end
      12'b000111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_449;
      end
      12'b000111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_450;
      end
      12'b000111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_451;
      end
      12'b000111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_452;
      end
      12'b000111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_453;
      end
      12'b000111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_454;
      end
      12'b000111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_455;
      end
      12'b000111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_456;
      end
      12'b000111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_457;
      end
      12'b000111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_458;
      end
      12'b000111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_459;
      end
      12'b000111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_460;
      end
      12'b000111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_461;
      end
      12'b000111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_462;
      end
      12'b000111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_463;
      end
      12'b000111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_464;
      end
      12'b000111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_465;
      end
      12'b000111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_466;
      end
      12'b000111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_467;
      end
      12'b000111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_468;
      end
      12'b000111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_469;
      end
      12'b000111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_470;
      end
      12'b000111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_471;
      end
      12'b000111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_472;
      end
      12'b000111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_473;
      end
      12'b000111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_474;
      end
      12'b000111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_475;
      end
      12'b000111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_476;
      end
      12'b000111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_477;
      end
      12'b000111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_478;
      end
      12'b000111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_479;
      end
      12'b000111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_480;
      end
      12'b000111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_481;
      end
      12'b000111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_482;
      end
      12'b000111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_483;
      end
      12'b000111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_484;
      end
      12'b000111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_485;
      end
      12'b000111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_486;
      end
      12'b000111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_487;
      end
      12'b000111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_488;
      end
      12'b000111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_489;
      end
      12'b000111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_490;
      end
      12'b000111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_491;
      end
      12'b000111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_492;
      end
      12'b000111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_493;
      end
      12'b000111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_494;
      end
      12'b000111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_495;
      end
      12'b000111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_496;
      end
      12'b000111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_497;
      end
      12'b000111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_498;
      end
      12'b000111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_499;
      end
      12'b000111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_500;
      end
      12'b000111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_501;
      end
      12'b000111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_502;
      end
      12'b000111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_503;
      end
      12'b000111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_504;
      end
      12'b000111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_505;
      end
      12'b000111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_506;
      end
      12'b000111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_507;
      end
      12'b000111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_508;
      end
      12'b000111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_509;
      end
      12'b000111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_510;
      end
      12'b000111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_511;
      end
      12'b001000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_512;
      end
      12'b001000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_513;
      end
      12'b001000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_514;
      end
      12'b001000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_515;
      end
      12'b001000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_516;
      end
      12'b001000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_517;
      end
      12'b001000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_518;
      end
      12'b001000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_519;
      end
      12'b001000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_520;
      end
      12'b001000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_521;
      end
      12'b001000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_522;
      end
      12'b001000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_523;
      end
      12'b001000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_524;
      end
      12'b001000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_525;
      end
      12'b001000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_526;
      end
      12'b001000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_527;
      end
      12'b001000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_528;
      end
      12'b001000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_529;
      end
      12'b001000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_530;
      end
      12'b001000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_531;
      end
      12'b001000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_532;
      end
      12'b001000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_533;
      end
      12'b001000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_534;
      end
      12'b001000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_535;
      end
      12'b001000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_536;
      end
      12'b001000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_537;
      end
      12'b001000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_538;
      end
      12'b001000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_539;
      end
      12'b001000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_540;
      end
      12'b001000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_541;
      end
      12'b001000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_542;
      end
      12'b001000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_543;
      end
      12'b001000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_544;
      end
      12'b001000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_545;
      end
      12'b001000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_546;
      end
      12'b001000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_547;
      end
      12'b001000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_548;
      end
      12'b001000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_549;
      end
      12'b001000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_550;
      end
      12'b001000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_551;
      end
      12'b001000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_552;
      end
      12'b001000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_553;
      end
      12'b001000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_554;
      end
      12'b001000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_555;
      end
      12'b001000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_556;
      end
      12'b001000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_557;
      end
      12'b001000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_558;
      end
      12'b001000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_559;
      end
      12'b001000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_560;
      end
      12'b001000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_561;
      end
      12'b001000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_562;
      end
      12'b001000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_563;
      end
      12'b001000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_564;
      end
      12'b001000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_565;
      end
      12'b001000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_566;
      end
      12'b001000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_567;
      end
      12'b001000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_568;
      end
      12'b001000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_569;
      end
      12'b001000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_570;
      end
      12'b001000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_571;
      end
      12'b001000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_572;
      end
      12'b001000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_573;
      end
      12'b001000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_574;
      end
      12'b001000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_575;
      end
      12'b001001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_576;
      end
      12'b001001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_577;
      end
      12'b001001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_578;
      end
      12'b001001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_579;
      end
      12'b001001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_580;
      end
      12'b001001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_581;
      end
      12'b001001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_582;
      end
      12'b001001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_583;
      end
      12'b001001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_584;
      end
      12'b001001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_585;
      end
      12'b001001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_586;
      end
      12'b001001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_587;
      end
      12'b001001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_588;
      end
      12'b001001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_589;
      end
      12'b001001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_590;
      end
      12'b001001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_591;
      end
      12'b001001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_592;
      end
      12'b001001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_593;
      end
      12'b001001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_594;
      end
      12'b001001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_595;
      end
      12'b001001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_596;
      end
      12'b001001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_597;
      end
      12'b001001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_598;
      end
      12'b001001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_599;
      end
      12'b001001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_600;
      end
      12'b001001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_601;
      end
      12'b001001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_602;
      end
      12'b001001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_603;
      end
      12'b001001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_604;
      end
      12'b001001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_605;
      end
      12'b001001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_606;
      end
      12'b001001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_607;
      end
      12'b001001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_608;
      end
      12'b001001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_609;
      end
      12'b001001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_610;
      end
      12'b001001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_611;
      end
      12'b001001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_612;
      end
      12'b001001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_613;
      end
      12'b001001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_614;
      end
      12'b001001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_615;
      end
      12'b001001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_616;
      end
      12'b001001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_617;
      end
      12'b001001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_618;
      end
      12'b001001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_619;
      end
      12'b001001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_620;
      end
      12'b001001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_621;
      end
      12'b001001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_622;
      end
      12'b001001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_623;
      end
      12'b001001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_624;
      end
      12'b001001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_625;
      end
      12'b001001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_626;
      end
      12'b001001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_627;
      end
      12'b001001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_628;
      end
      12'b001001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_629;
      end
      12'b001001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_630;
      end
      12'b001001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_631;
      end
      12'b001001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_632;
      end
      12'b001001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_633;
      end
      12'b001001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_634;
      end
      12'b001001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_635;
      end
      12'b001001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_636;
      end
      12'b001001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_637;
      end
      12'b001001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_638;
      end
      12'b001001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_639;
      end
      12'b001010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_640;
      end
      12'b001010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_641;
      end
      12'b001010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_642;
      end
      12'b001010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_643;
      end
      12'b001010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_644;
      end
      12'b001010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_645;
      end
      12'b001010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_646;
      end
      12'b001010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_647;
      end
      12'b001010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_648;
      end
      12'b001010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_649;
      end
      12'b001010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_650;
      end
      12'b001010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_651;
      end
      12'b001010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_652;
      end
      12'b001010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_653;
      end
      12'b001010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_654;
      end
      12'b001010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_655;
      end
      12'b001010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_656;
      end
      12'b001010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_657;
      end
      12'b001010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_658;
      end
      12'b001010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_659;
      end
      12'b001010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_660;
      end
      12'b001010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_661;
      end
      12'b001010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_662;
      end
      12'b001010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_663;
      end
      12'b001010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_664;
      end
      12'b001010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_665;
      end
      12'b001010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_666;
      end
      12'b001010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_667;
      end
      12'b001010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_668;
      end
      12'b001010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_669;
      end
      12'b001010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_670;
      end
      12'b001010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_671;
      end
      12'b001010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_672;
      end
      12'b001010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_673;
      end
      12'b001010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_674;
      end
      12'b001010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_675;
      end
      12'b001010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_676;
      end
      12'b001010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_677;
      end
      12'b001010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_678;
      end
      12'b001010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_679;
      end
      12'b001010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_680;
      end
      12'b001010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_681;
      end
      12'b001010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_682;
      end
      12'b001010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_683;
      end
      12'b001010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_684;
      end
      12'b001010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_685;
      end
      12'b001010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_686;
      end
      12'b001010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_687;
      end
      12'b001010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_688;
      end
      12'b001010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_689;
      end
      12'b001010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_690;
      end
      12'b001010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_691;
      end
      12'b001010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_692;
      end
      12'b001010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_693;
      end
      12'b001010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_694;
      end
      12'b001010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_695;
      end
      12'b001010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_696;
      end
      12'b001010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_697;
      end
      12'b001010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_698;
      end
      12'b001010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_699;
      end
      12'b001010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_700;
      end
      12'b001010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_701;
      end
      12'b001010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_702;
      end
      12'b001010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_703;
      end
      12'b001011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_704;
      end
      12'b001011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_705;
      end
      12'b001011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_706;
      end
      12'b001011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_707;
      end
      12'b001011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_708;
      end
      12'b001011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_709;
      end
      12'b001011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_710;
      end
      12'b001011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_711;
      end
      12'b001011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_712;
      end
      12'b001011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_713;
      end
      12'b001011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_714;
      end
      12'b001011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_715;
      end
      12'b001011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_716;
      end
      12'b001011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_717;
      end
      12'b001011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_718;
      end
      12'b001011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_719;
      end
      12'b001011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_720;
      end
      12'b001011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_721;
      end
      12'b001011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_722;
      end
      12'b001011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_723;
      end
      12'b001011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_724;
      end
      12'b001011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_725;
      end
      12'b001011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_726;
      end
      12'b001011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_727;
      end
      12'b001011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_728;
      end
      12'b001011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_729;
      end
      12'b001011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_730;
      end
      12'b001011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_731;
      end
      12'b001011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_732;
      end
      12'b001011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_733;
      end
      12'b001011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_734;
      end
      12'b001011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_735;
      end
      12'b001011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_736;
      end
      12'b001011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_737;
      end
      12'b001011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_738;
      end
      12'b001011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_739;
      end
      12'b001011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_740;
      end
      12'b001011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_741;
      end
      12'b001011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_742;
      end
      12'b001011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_743;
      end
      12'b001011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_744;
      end
      12'b001011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_745;
      end
      12'b001011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_746;
      end
      12'b001011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_747;
      end
      12'b001011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_748;
      end
      12'b001011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_749;
      end
      12'b001011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_750;
      end
      12'b001011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_751;
      end
      12'b001011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_752;
      end
      12'b001011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_753;
      end
      12'b001011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_754;
      end
      12'b001011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_755;
      end
      12'b001011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_756;
      end
      12'b001011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_757;
      end
      12'b001011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_758;
      end
      12'b001011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_759;
      end
      12'b001011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_760;
      end
      12'b001011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_761;
      end
      12'b001011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_762;
      end
      12'b001011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_763;
      end
      12'b001011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_764;
      end
      12'b001011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_765;
      end
      12'b001011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_766;
      end
      12'b001011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_767;
      end
      12'b001100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_768;
      end
      12'b001100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_769;
      end
      12'b001100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_770;
      end
      12'b001100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_771;
      end
      12'b001100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_772;
      end
      12'b001100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_773;
      end
      12'b001100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_774;
      end
      12'b001100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_775;
      end
      12'b001100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_776;
      end
      12'b001100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_777;
      end
      12'b001100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_778;
      end
      12'b001100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_779;
      end
      12'b001100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_780;
      end
      12'b001100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_781;
      end
      12'b001100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_782;
      end
      12'b001100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_783;
      end
      12'b001100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_784;
      end
      12'b001100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_785;
      end
      12'b001100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_786;
      end
      12'b001100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_787;
      end
      12'b001100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_788;
      end
      12'b001100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_789;
      end
      12'b001100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_790;
      end
      12'b001100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_791;
      end
      12'b001100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_792;
      end
      12'b001100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_793;
      end
      12'b001100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_794;
      end
      12'b001100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_795;
      end
      12'b001100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_796;
      end
      12'b001100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_797;
      end
      12'b001100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_798;
      end
      12'b001100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_799;
      end
      12'b001100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_800;
      end
      12'b001100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_801;
      end
      12'b001100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_802;
      end
      12'b001100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_803;
      end
      12'b001100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_804;
      end
      12'b001100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_805;
      end
      12'b001100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_806;
      end
      12'b001100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_807;
      end
      12'b001100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_808;
      end
      12'b001100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_809;
      end
      12'b001100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_810;
      end
      12'b001100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_811;
      end
      12'b001100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_812;
      end
      12'b001100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_813;
      end
      12'b001100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_814;
      end
      12'b001100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_815;
      end
      12'b001100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_816;
      end
      12'b001100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_817;
      end
      12'b001100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_818;
      end
      12'b001100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_819;
      end
      12'b001100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_820;
      end
      12'b001100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_821;
      end
      12'b001100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_822;
      end
      12'b001100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_823;
      end
      12'b001100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_824;
      end
      12'b001100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_825;
      end
      12'b001100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_826;
      end
      12'b001100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_827;
      end
      12'b001100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_828;
      end
      12'b001100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_829;
      end
      12'b001100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_830;
      end
      12'b001100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_831;
      end
      12'b001101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_832;
      end
      12'b001101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_833;
      end
      12'b001101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_834;
      end
      12'b001101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_835;
      end
      12'b001101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_836;
      end
      12'b001101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_837;
      end
      12'b001101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_838;
      end
      12'b001101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_839;
      end
      12'b001101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_840;
      end
      12'b001101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_841;
      end
      12'b001101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_842;
      end
      12'b001101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_843;
      end
      12'b001101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_844;
      end
      12'b001101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_845;
      end
      12'b001101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_846;
      end
      12'b001101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_847;
      end
      12'b001101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_848;
      end
      12'b001101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_849;
      end
      12'b001101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_850;
      end
      12'b001101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_851;
      end
      12'b001101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_852;
      end
      12'b001101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_853;
      end
      12'b001101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_854;
      end
      12'b001101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_855;
      end
      12'b001101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_856;
      end
      12'b001101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_857;
      end
      12'b001101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_858;
      end
      12'b001101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_859;
      end
      12'b001101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_860;
      end
      12'b001101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_861;
      end
      12'b001101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_862;
      end
      12'b001101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_863;
      end
      12'b001101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_864;
      end
      12'b001101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_865;
      end
      12'b001101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_866;
      end
      12'b001101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_867;
      end
      12'b001101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_868;
      end
      12'b001101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_869;
      end
      12'b001101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_870;
      end
      12'b001101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_871;
      end
      12'b001101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_872;
      end
      12'b001101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_873;
      end
      12'b001101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_874;
      end
      12'b001101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_875;
      end
      12'b001101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_876;
      end
      12'b001101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_877;
      end
      12'b001101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_878;
      end
      12'b001101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_879;
      end
      12'b001101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_880;
      end
      12'b001101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_881;
      end
      12'b001101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_882;
      end
      12'b001101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_883;
      end
      12'b001101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_884;
      end
      12'b001101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_885;
      end
      12'b001101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_886;
      end
      12'b001101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_887;
      end
      12'b001101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_888;
      end
      12'b001101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_889;
      end
      12'b001101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_890;
      end
      12'b001101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_891;
      end
      12'b001101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_892;
      end
      12'b001101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_893;
      end
      12'b001101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_894;
      end
      12'b001101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_895;
      end
      12'b001110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_896;
      end
      12'b001110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_897;
      end
      12'b001110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_898;
      end
      12'b001110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_899;
      end
      12'b001110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_900;
      end
      12'b001110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_901;
      end
      12'b001110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_902;
      end
      12'b001110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_903;
      end
      12'b001110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_904;
      end
      12'b001110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_905;
      end
      12'b001110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_906;
      end
      12'b001110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_907;
      end
      12'b001110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_908;
      end
      12'b001110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_909;
      end
      12'b001110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_910;
      end
      12'b001110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_911;
      end
      12'b001110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_912;
      end
      12'b001110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_913;
      end
      12'b001110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_914;
      end
      12'b001110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_915;
      end
      12'b001110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_916;
      end
      12'b001110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_917;
      end
      12'b001110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_918;
      end
      12'b001110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_919;
      end
      12'b001110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_920;
      end
      12'b001110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_921;
      end
      12'b001110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_922;
      end
      12'b001110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_923;
      end
      12'b001110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_924;
      end
      12'b001110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_925;
      end
      12'b001110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_926;
      end
      12'b001110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_927;
      end
      12'b001110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_928;
      end
      12'b001110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_929;
      end
      12'b001110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_930;
      end
      12'b001110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_931;
      end
      12'b001110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_932;
      end
      12'b001110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_933;
      end
      12'b001110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_934;
      end
      12'b001110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_935;
      end
      12'b001110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_936;
      end
      12'b001110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_937;
      end
      12'b001110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_938;
      end
      12'b001110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_939;
      end
      12'b001110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_940;
      end
      12'b001110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_941;
      end
      12'b001110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_942;
      end
      12'b001110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_943;
      end
      12'b001110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_944;
      end
      12'b001110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_945;
      end
      12'b001110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_946;
      end
      12'b001110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_947;
      end
      12'b001110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_948;
      end
      12'b001110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_949;
      end
      12'b001110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_950;
      end
      12'b001110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_951;
      end
      12'b001110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_952;
      end
      12'b001110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_953;
      end
      12'b001110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_954;
      end
      12'b001110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_955;
      end
      12'b001110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_956;
      end
      12'b001110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_957;
      end
      12'b001110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_958;
      end
      12'b001110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_959;
      end
      12'b001111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_960;
      end
      12'b001111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_961;
      end
      12'b001111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_962;
      end
      12'b001111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_963;
      end
      12'b001111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_964;
      end
      12'b001111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_965;
      end
      12'b001111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_966;
      end
      12'b001111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_967;
      end
      12'b001111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_968;
      end
      12'b001111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_969;
      end
      12'b001111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_970;
      end
      12'b001111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_971;
      end
      12'b001111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_972;
      end
      12'b001111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_973;
      end
      12'b001111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_974;
      end
      12'b001111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_975;
      end
      12'b001111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_976;
      end
      12'b001111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_977;
      end
      12'b001111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_978;
      end
      12'b001111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_979;
      end
      12'b001111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_980;
      end
      12'b001111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_981;
      end
      12'b001111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_982;
      end
      12'b001111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_983;
      end
      12'b001111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_984;
      end
      12'b001111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_985;
      end
      12'b001111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_986;
      end
      12'b001111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_987;
      end
      12'b001111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_988;
      end
      12'b001111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_989;
      end
      12'b001111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_990;
      end
      12'b001111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_991;
      end
      12'b001111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_992;
      end
      12'b001111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_993;
      end
      12'b001111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_994;
      end
      12'b001111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_995;
      end
      12'b001111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_996;
      end
      12'b001111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_997;
      end
      12'b001111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_998;
      end
      12'b001111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_999;
      end
      12'b001111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1000;
      end
      12'b001111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1001;
      end
      12'b001111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1002;
      end
      12'b001111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1003;
      end
      12'b001111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1004;
      end
      12'b001111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1005;
      end
      12'b001111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1006;
      end
      12'b001111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1007;
      end
      12'b001111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1008;
      end
      12'b001111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1009;
      end
      12'b001111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1010;
      end
      12'b001111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1011;
      end
      12'b001111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1012;
      end
      12'b001111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1013;
      end
      12'b001111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1014;
      end
      12'b001111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1015;
      end
      12'b001111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1016;
      end
      12'b001111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1017;
      end
      12'b001111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1018;
      end
      12'b001111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1019;
      end
      12'b001111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1020;
      end
      12'b001111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1021;
      end
      12'b001111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1022;
      end
      12'b001111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1023;
      end
      12'b010000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1024;
      end
      12'b010000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1025;
      end
      12'b010000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1026;
      end
      12'b010000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1027;
      end
      12'b010000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1028;
      end
      12'b010000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1029;
      end
      12'b010000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1030;
      end
      12'b010000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1031;
      end
      12'b010000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1032;
      end
      12'b010000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1033;
      end
      12'b010000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1034;
      end
      12'b010000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1035;
      end
      12'b010000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1036;
      end
      12'b010000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1037;
      end
      12'b010000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1038;
      end
      12'b010000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1039;
      end
      12'b010000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1040;
      end
      12'b010000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1041;
      end
      12'b010000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1042;
      end
      12'b010000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1043;
      end
      12'b010000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1044;
      end
      12'b010000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1045;
      end
      12'b010000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1046;
      end
      12'b010000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1047;
      end
      12'b010000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1048;
      end
      12'b010000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1049;
      end
      12'b010000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1050;
      end
      12'b010000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1051;
      end
      12'b010000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1052;
      end
      12'b010000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1053;
      end
      12'b010000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1054;
      end
      12'b010000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1055;
      end
      12'b010000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1056;
      end
      12'b010000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1057;
      end
      12'b010000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1058;
      end
      12'b010000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1059;
      end
      12'b010000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1060;
      end
      12'b010000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1061;
      end
      12'b010000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1062;
      end
      12'b010000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1063;
      end
      12'b010000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1064;
      end
      12'b010000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1065;
      end
      12'b010000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1066;
      end
      12'b010000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1067;
      end
      12'b010000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1068;
      end
      12'b010000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1069;
      end
      12'b010000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1070;
      end
      12'b010000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1071;
      end
      12'b010000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1072;
      end
      12'b010000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1073;
      end
      12'b010000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1074;
      end
      12'b010000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1075;
      end
      12'b010000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1076;
      end
      12'b010000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1077;
      end
      12'b010000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1078;
      end
      12'b010000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1079;
      end
      12'b010000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1080;
      end
      12'b010000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1081;
      end
      12'b010000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1082;
      end
      12'b010000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1083;
      end
      12'b010000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1084;
      end
      12'b010000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1085;
      end
      12'b010000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1086;
      end
      12'b010000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1087;
      end
      12'b010001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1088;
      end
      12'b010001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1089;
      end
      12'b010001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1090;
      end
      12'b010001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1091;
      end
      12'b010001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1092;
      end
      12'b010001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1093;
      end
      12'b010001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1094;
      end
      12'b010001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1095;
      end
      12'b010001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1096;
      end
      12'b010001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1097;
      end
      12'b010001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1098;
      end
      12'b010001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1099;
      end
      12'b010001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1100;
      end
      12'b010001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1101;
      end
      12'b010001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1102;
      end
      12'b010001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1103;
      end
      12'b010001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1104;
      end
      12'b010001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1105;
      end
      12'b010001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1106;
      end
      12'b010001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1107;
      end
      12'b010001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1108;
      end
      12'b010001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1109;
      end
      12'b010001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1110;
      end
      12'b010001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1111;
      end
      12'b010001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1112;
      end
      12'b010001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1113;
      end
      12'b010001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1114;
      end
      12'b010001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1115;
      end
      12'b010001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1116;
      end
      12'b010001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1117;
      end
      12'b010001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1118;
      end
      12'b010001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1119;
      end
      12'b010001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1120;
      end
      12'b010001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1121;
      end
      12'b010001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1122;
      end
      12'b010001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1123;
      end
      12'b010001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1124;
      end
      12'b010001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1125;
      end
      12'b010001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1126;
      end
      12'b010001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1127;
      end
      12'b010001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1128;
      end
      12'b010001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1129;
      end
      12'b010001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1130;
      end
      12'b010001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1131;
      end
      12'b010001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1132;
      end
      12'b010001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1133;
      end
      12'b010001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1134;
      end
      12'b010001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1135;
      end
      12'b010001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1136;
      end
      12'b010001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1137;
      end
      12'b010001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1138;
      end
      12'b010001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1139;
      end
      12'b010001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1140;
      end
      12'b010001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1141;
      end
      12'b010001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1142;
      end
      12'b010001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1143;
      end
      12'b010001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1144;
      end
      12'b010001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1145;
      end
      12'b010001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1146;
      end
      12'b010001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1147;
      end
      12'b010001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1148;
      end
      12'b010001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1149;
      end
      12'b010001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1150;
      end
      12'b010001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1151;
      end
      12'b010010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1152;
      end
      12'b010010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1153;
      end
      12'b010010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1154;
      end
      12'b010010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1155;
      end
      12'b010010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1156;
      end
      12'b010010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1157;
      end
      12'b010010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1158;
      end
      12'b010010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1159;
      end
      12'b010010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1160;
      end
      12'b010010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1161;
      end
      12'b010010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1162;
      end
      12'b010010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1163;
      end
      12'b010010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1164;
      end
      12'b010010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1165;
      end
      12'b010010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1166;
      end
      12'b010010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1167;
      end
      12'b010010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1168;
      end
      12'b010010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1169;
      end
      12'b010010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1170;
      end
      12'b010010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1171;
      end
      12'b010010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1172;
      end
      12'b010010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1173;
      end
      12'b010010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1174;
      end
      12'b010010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1175;
      end
      12'b010010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1176;
      end
      12'b010010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1177;
      end
      12'b010010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1178;
      end
      12'b010010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1179;
      end
      12'b010010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1180;
      end
      12'b010010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1181;
      end
      12'b010010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1182;
      end
      12'b010010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1183;
      end
      12'b010010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1184;
      end
      12'b010010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1185;
      end
      12'b010010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1186;
      end
      12'b010010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1187;
      end
      12'b010010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1188;
      end
      12'b010010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1189;
      end
      12'b010010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1190;
      end
      12'b010010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1191;
      end
      12'b010010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1192;
      end
      12'b010010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1193;
      end
      12'b010010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1194;
      end
      12'b010010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1195;
      end
      12'b010010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1196;
      end
      12'b010010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1197;
      end
      12'b010010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1198;
      end
      12'b010010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1199;
      end
      12'b010010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1200;
      end
      12'b010010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1201;
      end
      12'b010010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1202;
      end
      12'b010010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1203;
      end
      12'b010010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1204;
      end
      12'b010010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1205;
      end
      12'b010010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1206;
      end
      12'b010010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1207;
      end
      12'b010010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1208;
      end
      12'b010010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1209;
      end
      12'b010010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1210;
      end
      12'b010010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1211;
      end
      12'b010010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1212;
      end
      12'b010010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1213;
      end
      12'b010010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1214;
      end
      12'b010010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1215;
      end
      12'b010011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1216;
      end
      12'b010011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1217;
      end
      12'b010011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1218;
      end
      12'b010011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1219;
      end
      12'b010011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1220;
      end
      12'b010011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1221;
      end
      12'b010011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1222;
      end
      12'b010011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1223;
      end
      12'b010011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1224;
      end
      12'b010011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1225;
      end
      12'b010011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1226;
      end
      12'b010011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1227;
      end
      12'b010011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1228;
      end
      12'b010011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1229;
      end
      12'b010011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1230;
      end
      12'b010011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1231;
      end
      12'b010011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1232;
      end
      12'b010011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1233;
      end
      12'b010011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1234;
      end
      12'b010011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1235;
      end
      12'b010011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1236;
      end
      12'b010011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1237;
      end
      12'b010011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1238;
      end
      12'b010011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1239;
      end
      12'b010011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1240;
      end
      12'b010011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1241;
      end
      12'b010011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1242;
      end
      12'b010011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1243;
      end
      12'b010011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1244;
      end
      12'b010011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1245;
      end
      12'b010011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1246;
      end
      12'b010011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1247;
      end
      12'b010011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1248;
      end
      12'b010011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1249;
      end
      12'b010011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1250;
      end
      12'b010011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1251;
      end
      12'b010011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1252;
      end
      12'b010011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1253;
      end
      12'b010011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1254;
      end
      12'b010011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1255;
      end
      12'b010011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1256;
      end
      12'b010011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1257;
      end
      12'b010011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1258;
      end
      12'b010011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1259;
      end
      12'b010011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1260;
      end
      12'b010011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1261;
      end
      12'b010011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1262;
      end
      12'b010011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1263;
      end
      12'b010011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1264;
      end
      12'b010011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1265;
      end
      12'b010011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1266;
      end
      12'b010011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1267;
      end
      12'b010011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1268;
      end
      12'b010011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1269;
      end
      12'b010011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1270;
      end
      12'b010011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1271;
      end
      12'b010011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1272;
      end
      12'b010011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1273;
      end
      12'b010011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1274;
      end
      12'b010011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1275;
      end
      12'b010011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1276;
      end
      12'b010011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1277;
      end
      12'b010011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1278;
      end
      12'b010011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1279;
      end
      12'b010100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1280;
      end
      12'b010100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1281;
      end
      12'b010100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1282;
      end
      12'b010100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1283;
      end
      12'b010100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1284;
      end
      12'b010100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1285;
      end
      12'b010100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1286;
      end
      12'b010100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1287;
      end
      12'b010100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1288;
      end
      12'b010100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1289;
      end
      12'b010100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1290;
      end
      12'b010100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1291;
      end
      12'b010100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1292;
      end
      12'b010100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1293;
      end
      12'b010100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1294;
      end
      12'b010100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1295;
      end
      12'b010100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1296;
      end
      12'b010100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1297;
      end
      12'b010100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1298;
      end
      12'b010100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1299;
      end
      12'b010100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1300;
      end
      12'b010100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1301;
      end
      12'b010100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1302;
      end
      12'b010100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1303;
      end
      12'b010100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1304;
      end
      12'b010100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1305;
      end
      12'b010100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1306;
      end
      12'b010100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1307;
      end
      12'b010100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1308;
      end
      12'b010100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1309;
      end
      12'b010100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1310;
      end
      12'b010100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1311;
      end
      12'b010100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1312;
      end
      12'b010100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1313;
      end
      12'b010100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1314;
      end
      12'b010100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1315;
      end
      12'b010100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1316;
      end
      12'b010100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1317;
      end
      12'b010100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1318;
      end
      12'b010100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1319;
      end
      12'b010100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1320;
      end
      12'b010100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1321;
      end
      12'b010100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1322;
      end
      12'b010100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1323;
      end
      12'b010100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1324;
      end
      12'b010100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1325;
      end
      12'b010100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1326;
      end
      12'b010100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1327;
      end
      12'b010100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1328;
      end
      12'b010100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1329;
      end
      12'b010100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1330;
      end
      12'b010100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1331;
      end
      12'b010100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1332;
      end
      12'b010100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1333;
      end
      12'b010100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1334;
      end
      12'b010100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1335;
      end
      12'b010100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1336;
      end
      12'b010100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1337;
      end
      12'b010100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1338;
      end
      12'b010100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1339;
      end
      12'b010100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1340;
      end
      12'b010100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1341;
      end
      12'b010100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1342;
      end
      12'b010100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1343;
      end
      12'b010101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1344;
      end
      12'b010101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1345;
      end
      12'b010101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1346;
      end
      12'b010101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1347;
      end
      12'b010101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1348;
      end
      12'b010101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1349;
      end
      12'b010101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1350;
      end
      12'b010101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1351;
      end
      12'b010101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1352;
      end
      12'b010101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1353;
      end
      12'b010101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1354;
      end
      12'b010101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1355;
      end
      12'b010101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1356;
      end
      12'b010101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1357;
      end
      12'b010101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1358;
      end
      12'b010101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1359;
      end
      12'b010101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1360;
      end
      12'b010101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1361;
      end
      12'b010101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1362;
      end
      12'b010101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1363;
      end
      12'b010101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1364;
      end
      12'b010101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1365;
      end
      12'b010101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1366;
      end
      12'b010101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1367;
      end
      12'b010101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1368;
      end
      12'b010101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1369;
      end
      12'b010101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1370;
      end
      12'b010101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1371;
      end
      12'b010101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1372;
      end
      12'b010101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1373;
      end
      12'b010101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1374;
      end
      12'b010101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1375;
      end
      12'b010101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1376;
      end
      12'b010101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1377;
      end
      12'b010101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1378;
      end
      12'b010101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1379;
      end
      12'b010101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1380;
      end
      12'b010101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1381;
      end
      12'b010101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1382;
      end
      12'b010101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1383;
      end
      12'b010101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1384;
      end
      12'b010101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1385;
      end
      12'b010101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1386;
      end
      12'b010101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1387;
      end
      12'b010101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1388;
      end
      12'b010101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1389;
      end
      12'b010101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1390;
      end
      12'b010101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1391;
      end
      12'b010101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1392;
      end
      12'b010101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1393;
      end
      12'b010101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1394;
      end
      12'b010101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1395;
      end
      12'b010101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1396;
      end
      12'b010101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1397;
      end
      12'b010101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1398;
      end
      12'b010101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1399;
      end
      12'b010101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1400;
      end
      12'b010101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1401;
      end
      12'b010101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1402;
      end
      12'b010101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1403;
      end
      12'b010101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1404;
      end
      12'b010101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1405;
      end
      12'b010101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1406;
      end
      12'b010101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1407;
      end
      12'b010110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1408;
      end
      12'b010110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1409;
      end
      12'b010110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1410;
      end
      12'b010110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1411;
      end
      12'b010110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1412;
      end
      12'b010110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1413;
      end
      12'b010110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1414;
      end
      12'b010110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1415;
      end
      12'b010110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1416;
      end
      12'b010110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1417;
      end
      12'b010110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1418;
      end
      12'b010110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1419;
      end
      12'b010110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1420;
      end
      12'b010110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1421;
      end
      12'b010110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1422;
      end
      12'b010110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1423;
      end
      12'b010110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1424;
      end
      12'b010110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1425;
      end
      12'b010110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1426;
      end
      12'b010110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1427;
      end
      12'b010110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1428;
      end
      12'b010110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1429;
      end
      12'b010110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1430;
      end
      12'b010110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1431;
      end
      12'b010110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1432;
      end
      12'b010110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1433;
      end
      12'b010110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1434;
      end
      12'b010110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1435;
      end
      12'b010110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1436;
      end
      12'b010110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1437;
      end
      12'b010110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1438;
      end
      12'b010110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1439;
      end
      12'b010110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1440;
      end
      12'b010110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1441;
      end
      12'b010110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1442;
      end
      12'b010110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1443;
      end
      12'b010110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1444;
      end
      12'b010110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1445;
      end
      12'b010110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1446;
      end
      12'b010110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1447;
      end
      12'b010110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1448;
      end
      12'b010110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1449;
      end
      12'b010110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1450;
      end
      12'b010110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1451;
      end
      12'b010110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1452;
      end
      12'b010110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1453;
      end
      12'b010110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1454;
      end
      12'b010110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1455;
      end
      12'b010110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1456;
      end
      12'b010110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1457;
      end
      12'b010110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1458;
      end
      12'b010110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1459;
      end
      12'b010110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1460;
      end
      12'b010110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1461;
      end
      12'b010110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1462;
      end
      12'b010110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1463;
      end
      12'b010110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1464;
      end
      12'b010110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1465;
      end
      12'b010110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1466;
      end
      12'b010110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1467;
      end
      12'b010110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1468;
      end
      12'b010110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1469;
      end
      12'b010110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1470;
      end
      12'b010110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1471;
      end
      12'b010111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1472;
      end
      12'b010111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1473;
      end
      12'b010111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1474;
      end
      12'b010111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1475;
      end
      12'b010111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1476;
      end
      12'b010111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1477;
      end
      12'b010111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1478;
      end
      12'b010111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1479;
      end
      12'b010111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1480;
      end
      12'b010111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1481;
      end
      12'b010111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1482;
      end
      12'b010111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1483;
      end
      12'b010111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1484;
      end
      12'b010111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1485;
      end
      12'b010111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1486;
      end
      12'b010111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1487;
      end
      12'b010111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1488;
      end
      12'b010111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1489;
      end
      12'b010111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1490;
      end
      12'b010111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1491;
      end
      12'b010111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1492;
      end
      12'b010111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1493;
      end
      12'b010111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1494;
      end
      12'b010111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1495;
      end
      12'b010111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1496;
      end
      12'b010111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1497;
      end
      12'b010111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1498;
      end
      12'b010111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1499;
      end
      12'b010111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1500;
      end
      12'b010111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1501;
      end
      12'b010111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1502;
      end
      12'b010111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1503;
      end
      12'b010111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1504;
      end
      12'b010111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1505;
      end
      12'b010111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1506;
      end
      12'b010111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1507;
      end
      12'b010111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1508;
      end
      12'b010111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1509;
      end
      12'b010111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1510;
      end
      12'b010111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1511;
      end
      12'b010111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1512;
      end
      12'b010111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1513;
      end
      12'b010111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1514;
      end
      12'b010111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1515;
      end
      12'b010111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1516;
      end
      12'b010111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1517;
      end
      12'b010111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1518;
      end
      12'b010111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1519;
      end
      12'b010111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1520;
      end
      12'b010111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1521;
      end
      12'b010111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1522;
      end
      12'b010111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1523;
      end
      12'b010111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1524;
      end
      12'b010111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1525;
      end
      12'b010111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1526;
      end
      12'b010111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1527;
      end
      12'b010111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1528;
      end
      12'b010111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1529;
      end
      12'b010111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1530;
      end
      12'b010111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1531;
      end
      12'b010111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1532;
      end
      12'b010111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1533;
      end
      12'b010111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1534;
      end
      12'b010111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1535;
      end
      12'b011000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1536;
      end
      12'b011000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1537;
      end
      12'b011000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1538;
      end
      12'b011000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1539;
      end
      12'b011000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1540;
      end
      12'b011000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1541;
      end
      12'b011000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1542;
      end
      12'b011000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1543;
      end
      12'b011000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1544;
      end
      12'b011000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1545;
      end
      12'b011000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1546;
      end
      12'b011000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1547;
      end
      12'b011000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1548;
      end
      12'b011000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1549;
      end
      12'b011000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1550;
      end
      12'b011000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1551;
      end
      12'b011000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1552;
      end
      12'b011000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1553;
      end
      12'b011000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1554;
      end
      12'b011000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1555;
      end
      12'b011000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1556;
      end
      12'b011000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1557;
      end
      12'b011000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1558;
      end
      12'b011000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1559;
      end
      12'b011000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1560;
      end
      12'b011000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1561;
      end
      12'b011000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1562;
      end
      12'b011000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1563;
      end
      12'b011000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1564;
      end
      12'b011000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1565;
      end
      12'b011000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1566;
      end
      12'b011000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1567;
      end
      12'b011000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1568;
      end
      12'b011000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1569;
      end
      12'b011000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1570;
      end
      12'b011000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1571;
      end
      12'b011000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1572;
      end
      12'b011000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1573;
      end
      12'b011000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1574;
      end
      12'b011000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1575;
      end
      12'b011000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1576;
      end
      12'b011000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1577;
      end
      12'b011000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1578;
      end
      12'b011000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1579;
      end
      12'b011000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1580;
      end
      12'b011000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1581;
      end
      12'b011000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1582;
      end
      12'b011000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1583;
      end
      12'b011000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1584;
      end
      12'b011000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1585;
      end
      12'b011000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1586;
      end
      12'b011000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1587;
      end
      12'b011000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1588;
      end
      12'b011000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1589;
      end
      12'b011000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1590;
      end
      12'b011000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1591;
      end
      12'b011000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1592;
      end
      12'b011000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1593;
      end
      12'b011000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1594;
      end
      12'b011000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1595;
      end
      12'b011000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1596;
      end
      12'b011000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1597;
      end
      12'b011000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1598;
      end
      12'b011000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1599;
      end
      12'b011001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1600;
      end
      12'b011001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1601;
      end
      12'b011001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1602;
      end
      12'b011001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1603;
      end
      12'b011001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1604;
      end
      12'b011001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1605;
      end
      12'b011001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1606;
      end
      12'b011001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1607;
      end
      12'b011001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1608;
      end
      12'b011001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1609;
      end
      12'b011001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1610;
      end
      12'b011001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1611;
      end
      12'b011001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1612;
      end
      12'b011001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1613;
      end
      12'b011001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1614;
      end
      12'b011001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1615;
      end
      12'b011001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1616;
      end
      12'b011001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1617;
      end
      12'b011001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1618;
      end
      12'b011001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1619;
      end
      12'b011001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1620;
      end
      12'b011001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1621;
      end
      12'b011001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1622;
      end
      12'b011001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1623;
      end
      12'b011001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1624;
      end
      12'b011001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1625;
      end
      12'b011001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1626;
      end
      12'b011001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1627;
      end
      12'b011001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1628;
      end
      12'b011001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1629;
      end
      12'b011001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1630;
      end
      12'b011001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1631;
      end
      12'b011001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1632;
      end
      12'b011001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1633;
      end
      12'b011001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1634;
      end
      12'b011001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1635;
      end
      12'b011001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1636;
      end
      12'b011001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1637;
      end
      12'b011001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1638;
      end
      12'b011001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1639;
      end
      12'b011001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1640;
      end
      12'b011001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1641;
      end
      12'b011001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1642;
      end
      12'b011001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1643;
      end
      12'b011001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1644;
      end
      12'b011001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1645;
      end
      12'b011001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1646;
      end
      12'b011001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1647;
      end
      12'b011001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1648;
      end
      12'b011001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1649;
      end
      12'b011001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1650;
      end
      12'b011001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1651;
      end
      12'b011001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1652;
      end
      12'b011001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1653;
      end
      12'b011001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1654;
      end
      12'b011001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1655;
      end
      12'b011001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1656;
      end
      12'b011001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1657;
      end
      12'b011001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1658;
      end
      12'b011001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1659;
      end
      12'b011001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1660;
      end
      12'b011001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1661;
      end
      12'b011001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1662;
      end
      12'b011001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1663;
      end
      12'b011010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1664;
      end
      12'b011010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1665;
      end
      12'b011010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1666;
      end
      12'b011010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1667;
      end
      12'b011010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1668;
      end
      12'b011010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1669;
      end
      12'b011010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1670;
      end
      12'b011010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1671;
      end
      12'b011010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1672;
      end
      12'b011010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1673;
      end
      12'b011010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1674;
      end
      12'b011010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1675;
      end
      12'b011010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1676;
      end
      12'b011010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1677;
      end
      12'b011010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1678;
      end
      12'b011010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1679;
      end
      12'b011010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1680;
      end
      12'b011010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1681;
      end
      12'b011010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1682;
      end
      12'b011010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1683;
      end
      12'b011010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1684;
      end
      12'b011010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1685;
      end
      12'b011010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1686;
      end
      12'b011010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1687;
      end
      12'b011010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1688;
      end
      12'b011010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1689;
      end
      12'b011010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1690;
      end
      12'b011010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1691;
      end
      12'b011010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1692;
      end
      12'b011010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1693;
      end
      12'b011010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1694;
      end
      12'b011010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1695;
      end
      12'b011010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1696;
      end
      12'b011010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1697;
      end
      12'b011010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1698;
      end
      12'b011010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1699;
      end
      12'b011010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1700;
      end
      12'b011010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1701;
      end
      12'b011010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1702;
      end
      12'b011010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1703;
      end
      12'b011010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1704;
      end
      12'b011010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1705;
      end
      12'b011010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1706;
      end
      12'b011010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1707;
      end
      12'b011010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1708;
      end
      12'b011010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1709;
      end
      12'b011010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1710;
      end
      12'b011010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1711;
      end
      12'b011010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1712;
      end
      12'b011010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1713;
      end
      12'b011010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1714;
      end
      12'b011010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1715;
      end
      12'b011010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1716;
      end
      12'b011010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1717;
      end
      12'b011010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1718;
      end
      12'b011010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1719;
      end
      12'b011010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1720;
      end
      12'b011010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1721;
      end
      12'b011010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1722;
      end
      12'b011010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1723;
      end
      12'b011010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1724;
      end
      12'b011010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1725;
      end
      12'b011010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1726;
      end
      12'b011010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1727;
      end
      12'b011011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1728;
      end
      12'b011011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1729;
      end
      12'b011011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1730;
      end
      12'b011011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1731;
      end
      12'b011011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1732;
      end
      12'b011011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1733;
      end
      12'b011011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1734;
      end
      12'b011011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1735;
      end
      12'b011011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1736;
      end
      12'b011011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1737;
      end
      12'b011011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1738;
      end
      12'b011011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1739;
      end
      12'b011011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1740;
      end
      12'b011011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1741;
      end
      12'b011011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1742;
      end
      12'b011011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1743;
      end
      12'b011011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1744;
      end
      12'b011011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1745;
      end
      12'b011011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1746;
      end
      12'b011011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1747;
      end
      12'b011011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1748;
      end
      12'b011011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1749;
      end
      12'b011011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1750;
      end
      12'b011011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1751;
      end
      12'b011011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1752;
      end
      12'b011011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1753;
      end
      12'b011011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1754;
      end
      12'b011011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1755;
      end
      12'b011011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1756;
      end
      12'b011011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1757;
      end
      12'b011011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1758;
      end
      12'b011011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1759;
      end
      12'b011011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1760;
      end
      12'b011011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1761;
      end
      12'b011011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1762;
      end
      12'b011011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1763;
      end
      12'b011011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1764;
      end
      12'b011011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1765;
      end
      12'b011011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1766;
      end
      12'b011011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1767;
      end
      12'b011011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1768;
      end
      12'b011011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1769;
      end
      12'b011011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1770;
      end
      12'b011011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1771;
      end
      12'b011011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1772;
      end
      12'b011011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1773;
      end
      12'b011011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1774;
      end
      12'b011011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1775;
      end
      12'b011011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1776;
      end
      12'b011011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1777;
      end
      12'b011011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1778;
      end
      12'b011011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1779;
      end
      12'b011011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1780;
      end
      12'b011011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1781;
      end
      12'b011011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1782;
      end
      12'b011011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1783;
      end
      12'b011011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1784;
      end
      12'b011011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1785;
      end
      12'b011011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1786;
      end
      12'b011011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1787;
      end
      12'b011011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1788;
      end
      12'b011011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1789;
      end
      12'b011011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1790;
      end
      12'b011011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1791;
      end
      12'b011100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1792;
      end
      12'b011100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1793;
      end
      12'b011100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1794;
      end
      12'b011100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1795;
      end
      12'b011100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1796;
      end
      12'b011100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1797;
      end
      12'b011100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1798;
      end
      12'b011100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1799;
      end
      12'b011100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1800;
      end
      12'b011100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1801;
      end
      12'b011100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1802;
      end
      12'b011100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1803;
      end
      12'b011100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1804;
      end
      12'b011100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1805;
      end
      12'b011100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1806;
      end
      12'b011100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1807;
      end
      12'b011100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1808;
      end
      12'b011100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1809;
      end
      12'b011100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1810;
      end
      12'b011100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1811;
      end
      12'b011100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1812;
      end
      12'b011100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1813;
      end
      12'b011100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1814;
      end
      12'b011100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1815;
      end
      12'b011100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1816;
      end
      12'b011100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1817;
      end
      12'b011100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1818;
      end
      12'b011100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1819;
      end
      12'b011100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1820;
      end
      12'b011100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1821;
      end
      12'b011100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1822;
      end
      12'b011100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1823;
      end
      12'b011100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1824;
      end
      12'b011100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1825;
      end
      12'b011100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1826;
      end
      12'b011100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1827;
      end
      12'b011100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1828;
      end
      12'b011100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1829;
      end
      12'b011100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1830;
      end
      12'b011100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1831;
      end
      12'b011100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1832;
      end
      12'b011100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1833;
      end
      12'b011100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1834;
      end
      12'b011100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1835;
      end
      12'b011100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1836;
      end
      12'b011100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1837;
      end
      12'b011100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1838;
      end
      12'b011100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1839;
      end
      12'b011100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1840;
      end
      12'b011100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1841;
      end
      12'b011100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1842;
      end
      12'b011100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1843;
      end
      12'b011100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1844;
      end
      12'b011100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1845;
      end
      12'b011100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1846;
      end
      12'b011100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1847;
      end
      12'b011100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1848;
      end
      12'b011100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1849;
      end
      12'b011100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1850;
      end
      12'b011100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1851;
      end
      12'b011100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1852;
      end
      12'b011100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1853;
      end
      12'b011100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1854;
      end
      12'b011100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1855;
      end
      12'b011101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1856;
      end
      12'b011101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1857;
      end
      12'b011101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1858;
      end
      12'b011101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1859;
      end
      12'b011101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1860;
      end
      12'b011101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1861;
      end
      12'b011101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1862;
      end
      12'b011101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1863;
      end
      12'b011101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1864;
      end
      12'b011101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1865;
      end
      12'b011101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1866;
      end
      12'b011101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1867;
      end
      12'b011101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1868;
      end
      12'b011101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1869;
      end
      12'b011101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1870;
      end
      12'b011101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1871;
      end
      12'b011101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1872;
      end
      12'b011101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1873;
      end
      12'b011101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1874;
      end
      12'b011101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1875;
      end
      12'b011101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1876;
      end
      12'b011101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1877;
      end
      12'b011101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1878;
      end
      12'b011101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1879;
      end
      12'b011101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1880;
      end
      12'b011101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1881;
      end
      12'b011101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1882;
      end
      12'b011101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1883;
      end
      12'b011101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1884;
      end
      12'b011101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1885;
      end
      12'b011101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1886;
      end
      12'b011101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1887;
      end
      12'b011101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1888;
      end
      12'b011101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1889;
      end
      12'b011101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1890;
      end
      12'b011101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1891;
      end
      12'b011101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1892;
      end
      12'b011101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1893;
      end
      12'b011101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1894;
      end
      12'b011101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1895;
      end
      12'b011101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1896;
      end
      12'b011101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1897;
      end
      12'b011101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1898;
      end
      12'b011101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1899;
      end
      12'b011101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1900;
      end
      12'b011101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1901;
      end
      12'b011101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1902;
      end
      12'b011101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1903;
      end
      12'b011101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1904;
      end
      12'b011101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1905;
      end
      12'b011101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1906;
      end
      12'b011101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1907;
      end
      12'b011101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1908;
      end
      12'b011101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1909;
      end
      12'b011101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1910;
      end
      12'b011101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1911;
      end
      12'b011101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1912;
      end
      12'b011101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1913;
      end
      12'b011101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1914;
      end
      12'b011101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1915;
      end
      12'b011101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1916;
      end
      12'b011101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1917;
      end
      12'b011101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1918;
      end
      12'b011101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1919;
      end
      12'b011110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1920;
      end
      12'b011110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1921;
      end
      12'b011110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1922;
      end
      12'b011110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1923;
      end
      12'b011110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1924;
      end
      12'b011110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1925;
      end
      12'b011110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1926;
      end
      12'b011110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1927;
      end
      12'b011110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1928;
      end
      12'b011110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1929;
      end
      12'b011110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1930;
      end
      12'b011110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1931;
      end
      12'b011110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1932;
      end
      12'b011110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1933;
      end
      12'b011110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1934;
      end
      12'b011110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1935;
      end
      12'b011110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1936;
      end
      12'b011110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1937;
      end
      12'b011110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1938;
      end
      12'b011110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1939;
      end
      12'b011110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1940;
      end
      12'b011110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1941;
      end
      12'b011110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1942;
      end
      12'b011110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1943;
      end
      12'b011110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1944;
      end
      12'b011110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1945;
      end
      12'b011110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1946;
      end
      12'b011110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1947;
      end
      12'b011110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1948;
      end
      12'b011110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1949;
      end
      12'b011110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1950;
      end
      12'b011110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1951;
      end
      12'b011110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1952;
      end
      12'b011110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1953;
      end
      12'b011110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1954;
      end
      12'b011110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1955;
      end
      12'b011110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1956;
      end
      12'b011110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1957;
      end
      12'b011110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1958;
      end
      12'b011110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1959;
      end
      12'b011110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1960;
      end
      12'b011110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1961;
      end
      12'b011110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1962;
      end
      12'b011110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1963;
      end
      12'b011110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1964;
      end
      12'b011110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1965;
      end
      12'b011110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1966;
      end
      12'b011110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1967;
      end
      12'b011110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1968;
      end
      12'b011110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1969;
      end
      12'b011110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1970;
      end
      12'b011110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1971;
      end
      12'b011110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1972;
      end
      12'b011110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1973;
      end
      12'b011110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1974;
      end
      12'b011110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1975;
      end
      12'b011110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1976;
      end
      12'b011110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1977;
      end
      12'b011110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1978;
      end
      12'b011110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1979;
      end
      12'b011110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1980;
      end
      12'b011110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1981;
      end
      12'b011110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1982;
      end
      12'b011110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1983;
      end
      12'b011111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1984;
      end
      12'b011111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1985;
      end
      12'b011111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1986;
      end
      12'b011111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1987;
      end
      12'b011111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1988;
      end
      12'b011111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1989;
      end
      12'b011111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1990;
      end
      12'b011111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1991;
      end
      12'b011111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_1992;
      end
      12'b011111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_1993;
      end
      12'b011111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_1994;
      end
      12'b011111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_1995;
      end
      12'b011111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_1996;
      end
      12'b011111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_1997;
      end
      12'b011111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_1998;
      end
      12'b011111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_1999;
      end
      12'b011111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2000;
      end
      12'b011111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2001;
      end
      12'b011111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2002;
      end
      12'b011111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2003;
      end
      12'b011111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2004;
      end
      12'b011111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2005;
      end
      12'b011111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2006;
      end
      12'b011111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2007;
      end
      12'b011111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2008;
      end
      12'b011111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2009;
      end
      12'b011111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2010;
      end
      12'b011111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2011;
      end
      12'b011111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2012;
      end
      12'b011111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2013;
      end
      12'b011111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2014;
      end
      12'b011111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2015;
      end
      12'b011111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2016;
      end
      12'b011111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2017;
      end
      12'b011111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2018;
      end
      12'b011111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2019;
      end
      12'b011111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2020;
      end
      12'b011111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2021;
      end
      12'b011111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2022;
      end
      12'b011111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2023;
      end
      12'b011111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2024;
      end
      12'b011111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2025;
      end
      12'b011111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2026;
      end
      12'b011111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2027;
      end
      12'b011111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2028;
      end
      12'b011111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2029;
      end
      12'b011111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2030;
      end
      12'b011111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2031;
      end
      12'b011111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2032;
      end
      12'b011111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2033;
      end
      12'b011111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2034;
      end
      12'b011111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2035;
      end
      12'b011111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2036;
      end
      12'b011111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2037;
      end
      12'b011111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2038;
      end
      12'b011111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2039;
      end
      12'b011111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2040;
      end
      12'b011111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2041;
      end
      12'b011111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2042;
      end
      12'b011111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2043;
      end
      12'b011111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2044;
      end
      12'b011111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2045;
      end
      12'b011111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2046;
      end
      12'b011111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2047;
      end
      12'b100000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2048;
      end
      12'b100000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2049;
      end
      12'b100000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2050;
      end
      12'b100000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2051;
      end
      12'b100000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2052;
      end
      12'b100000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2053;
      end
      12'b100000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2054;
      end
      12'b100000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2055;
      end
      12'b100000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2056;
      end
      12'b100000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2057;
      end
      12'b100000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2058;
      end
      12'b100000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2059;
      end
      12'b100000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2060;
      end
      12'b100000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2061;
      end
      12'b100000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2062;
      end
      12'b100000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2063;
      end
      12'b100000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2064;
      end
      12'b100000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2065;
      end
      12'b100000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2066;
      end
      12'b100000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2067;
      end
      12'b100000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2068;
      end
      12'b100000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2069;
      end
      12'b100000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2070;
      end
      12'b100000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2071;
      end
      12'b100000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2072;
      end
      12'b100000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2073;
      end
      12'b100000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2074;
      end
      12'b100000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2075;
      end
      12'b100000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2076;
      end
      12'b100000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2077;
      end
      12'b100000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2078;
      end
      12'b100000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2079;
      end
      12'b100000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2080;
      end
      12'b100000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2081;
      end
      12'b100000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2082;
      end
      12'b100000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2083;
      end
      12'b100000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2084;
      end
      12'b100000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2085;
      end
      12'b100000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2086;
      end
      12'b100000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2087;
      end
      12'b100000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2088;
      end
      12'b100000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2089;
      end
      12'b100000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2090;
      end
      12'b100000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2091;
      end
      12'b100000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2092;
      end
      12'b100000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2093;
      end
      12'b100000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2094;
      end
      12'b100000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2095;
      end
      12'b100000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2096;
      end
      12'b100000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2097;
      end
      12'b100000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2098;
      end
      12'b100000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2099;
      end
      12'b100000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2100;
      end
      12'b100000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2101;
      end
      12'b100000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2102;
      end
      12'b100000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2103;
      end
      12'b100000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2104;
      end
      12'b100000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2105;
      end
      12'b100000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2106;
      end
      12'b100000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2107;
      end
      12'b100000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2108;
      end
      12'b100000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2109;
      end
      12'b100000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2110;
      end
      12'b100000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2111;
      end
      12'b100001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2112;
      end
      12'b100001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2113;
      end
      12'b100001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2114;
      end
      12'b100001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2115;
      end
      12'b100001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2116;
      end
      12'b100001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2117;
      end
      12'b100001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2118;
      end
      12'b100001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2119;
      end
      12'b100001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2120;
      end
      12'b100001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2121;
      end
      12'b100001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2122;
      end
      12'b100001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2123;
      end
      12'b100001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2124;
      end
      12'b100001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2125;
      end
      12'b100001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2126;
      end
      12'b100001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2127;
      end
      12'b100001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2128;
      end
      12'b100001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2129;
      end
      12'b100001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2130;
      end
      12'b100001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2131;
      end
      12'b100001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2132;
      end
      12'b100001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2133;
      end
      12'b100001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2134;
      end
      12'b100001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2135;
      end
      12'b100001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2136;
      end
      12'b100001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2137;
      end
      12'b100001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2138;
      end
      12'b100001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2139;
      end
      12'b100001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2140;
      end
      12'b100001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2141;
      end
      12'b100001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2142;
      end
      12'b100001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2143;
      end
      12'b100001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2144;
      end
      12'b100001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2145;
      end
      12'b100001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2146;
      end
      12'b100001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2147;
      end
      12'b100001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2148;
      end
      12'b100001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2149;
      end
      12'b100001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2150;
      end
      12'b100001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2151;
      end
      12'b100001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2152;
      end
      12'b100001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2153;
      end
      12'b100001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2154;
      end
      12'b100001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2155;
      end
      12'b100001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2156;
      end
      12'b100001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2157;
      end
      12'b100001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2158;
      end
      12'b100001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2159;
      end
      12'b100001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2160;
      end
      12'b100001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2161;
      end
      12'b100001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2162;
      end
      12'b100001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2163;
      end
      12'b100001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2164;
      end
      12'b100001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2165;
      end
      12'b100001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2166;
      end
      12'b100001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2167;
      end
      12'b100001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2168;
      end
      12'b100001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2169;
      end
      12'b100001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2170;
      end
      12'b100001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2171;
      end
      12'b100001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2172;
      end
      12'b100001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2173;
      end
      12'b100001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2174;
      end
      12'b100001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2175;
      end
      12'b100010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2176;
      end
      12'b100010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2177;
      end
      12'b100010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2178;
      end
      12'b100010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2179;
      end
      12'b100010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2180;
      end
      12'b100010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2181;
      end
      12'b100010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2182;
      end
      12'b100010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2183;
      end
      12'b100010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2184;
      end
      12'b100010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2185;
      end
      12'b100010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2186;
      end
      12'b100010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2187;
      end
      12'b100010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2188;
      end
      12'b100010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2189;
      end
      12'b100010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2190;
      end
      12'b100010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2191;
      end
      12'b100010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2192;
      end
      12'b100010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2193;
      end
      12'b100010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2194;
      end
      12'b100010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2195;
      end
      12'b100010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2196;
      end
      12'b100010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2197;
      end
      12'b100010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2198;
      end
      12'b100010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2199;
      end
      12'b100010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2200;
      end
      12'b100010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2201;
      end
      12'b100010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2202;
      end
      12'b100010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2203;
      end
      12'b100010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2204;
      end
      12'b100010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2205;
      end
      12'b100010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2206;
      end
      12'b100010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2207;
      end
      12'b100010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2208;
      end
      12'b100010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2209;
      end
      12'b100010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2210;
      end
      12'b100010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2211;
      end
      12'b100010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2212;
      end
      12'b100010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2213;
      end
      12'b100010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2214;
      end
      12'b100010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2215;
      end
      12'b100010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2216;
      end
      12'b100010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2217;
      end
      12'b100010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2218;
      end
      12'b100010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2219;
      end
      12'b100010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2220;
      end
      12'b100010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2221;
      end
      12'b100010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2222;
      end
      12'b100010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2223;
      end
      12'b100010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2224;
      end
      12'b100010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2225;
      end
      12'b100010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2226;
      end
      12'b100010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2227;
      end
      12'b100010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2228;
      end
      12'b100010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2229;
      end
      12'b100010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2230;
      end
      12'b100010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2231;
      end
      12'b100010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2232;
      end
      12'b100010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2233;
      end
      12'b100010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2234;
      end
      12'b100010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2235;
      end
      12'b100010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2236;
      end
      12'b100010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2237;
      end
      12'b100010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2238;
      end
      12'b100010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2239;
      end
      12'b100011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2240;
      end
      12'b100011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2241;
      end
      12'b100011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2242;
      end
      12'b100011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2243;
      end
      12'b100011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2244;
      end
      12'b100011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2245;
      end
      12'b100011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2246;
      end
      12'b100011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2247;
      end
      12'b100011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2248;
      end
      12'b100011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2249;
      end
      12'b100011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2250;
      end
      12'b100011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2251;
      end
      12'b100011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2252;
      end
      12'b100011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2253;
      end
      12'b100011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2254;
      end
      12'b100011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2255;
      end
      12'b100011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2256;
      end
      12'b100011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2257;
      end
      12'b100011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2258;
      end
      12'b100011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2259;
      end
      12'b100011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2260;
      end
      12'b100011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2261;
      end
      12'b100011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2262;
      end
      12'b100011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2263;
      end
      12'b100011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2264;
      end
      12'b100011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2265;
      end
      12'b100011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2266;
      end
      12'b100011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2267;
      end
      12'b100011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2268;
      end
      12'b100011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2269;
      end
      12'b100011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2270;
      end
      12'b100011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2271;
      end
      12'b100011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2272;
      end
      12'b100011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2273;
      end
      12'b100011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2274;
      end
      12'b100011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2275;
      end
      12'b100011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2276;
      end
      12'b100011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2277;
      end
      12'b100011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2278;
      end
      12'b100011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2279;
      end
      12'b100011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2280;
      end
      12'b100011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2281;
      end
      12'b100011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2282;
      end
      12'b100011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2283;
      end
      12'b100011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2284;
      end
      12'b100011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2285;
      end
      12'b100011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2286;
      end
      12'b100011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2287;
      end
      12'b100011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2288;
      end
      12'b100011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2289;
      end
      12'b100011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2290;
      end
      12'b100011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2291;
      end
      12'b100011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2292;
      end
      12'b100011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2293;
      end
      12'b100011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2294;
      end
      12'b100011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2295;
      end
      12'b100011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2296;
      end
      12'b100011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2297;
      end
      12'b100011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2298;
      end
      12'b100011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2299;
      end
      12'b100011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2300;
      end
      12'b100011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2301;
      end
      12'b100011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2302;
      end
      12'b100011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2303;
      end
      12'b100100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2304;
      end
      12'b100100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2305;
      end
      12'b100100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2306;
      end
      12'b100100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2307;
      end
      12'b100100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2308;
      end
      12'b100100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2309;
      end
      12'b100100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2310;
      end
      12'b100100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2311;
      end
      12'b100100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2312;
      end
      12'b100100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2313;
      end
      12'b100100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2314;
      end
      12'b100100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2315;
      end
      12'b100100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2316;
      end
      12'b100100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2317;
      end
      12'b100100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2318;
      end
      12'b100100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2319;
      end
      12'b100100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2320;
      end
      12'b100100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2321;
      end
      12'b100100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2322;
      end
      12'b100100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2323;
      end
      12'b100100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2324;
      end
      12'b100100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2325;
      end
      12'b100100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2326;
      end
      12'b100100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2327;
      end
      12'b100100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2328;
      end
      12'b100100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2329;
      end
      12'b100100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2330;
      end
      12'b100100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2331;
      end
      12'b100100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2332;
      end
      12'b100100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2333;
      end
      12'b100100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2334;
      end
      12'b100100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2335;
      end
      12'b100100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2336;
      end
      12'b100100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2337;
      end
      12'b100100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2338;
      end
      12'b100100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2339;
      end
      12'b100100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2340;
      end
      12'b100100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2341;
      end
      12'b100100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2342;
      end
      12'b100100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2343;
      end
      12'b100100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2344;
      end
      12'b100100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2345;
      end
      12'b100100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2346;
      end
      12'b100100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2347;
      end
      12'b100100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2348;
      end
      12'b100100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2349;
      end
      12'b100100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2350;
      end
      12'b100100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2351;
      end
      12'b100100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2352;
      end
      12'b100100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2353;
      end
      12'b100100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2354;
      end
      12'b100100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2355;
      end
      12'b100100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2356;
      end
      12'b100100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2357;
      end
      12'b100100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2358;
      end
      12'b100100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2359;
      end
      12'b100100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2360;
      end
      12'b100100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2361;
      end
      12'b100100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2362;
      end
      12'b100100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2363;
      end
      12'b100100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2364;
      end
      12'b100100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2365;
      end
      12'b100100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2366;
      end
      12'b100100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2367;
      end
      12'b100101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2368;
      end
      12'b100101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2369;
      end
      12'b100101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2370;
      end
      12'b100101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2371;
      end
      12'b100101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2372;
      end
      12'b100101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2373;
      end
      12'b100101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2374;
      end
      12'b100101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2375;
      end
      12'b100101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2376;
      end
      12'b100101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2377;
      end
      12'b100101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2378;
      end
      12'b100101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2379;
      end
      12'b100101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2380;
      end
      12'b100101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2381;
      end
      12'b100101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2382;
      end
      12'b100101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2383;
      end
      12'b100101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2384;
      end
      12'b100101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2385;
      end
      12'b100101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2386;
      end
      12'b100101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2387;
      end
      12'b100101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2388;
      end
      12'b100101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2389;
      end
      12'b100101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2390;
      end
      12'b100101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2391;
      end
      12'b100101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2392;
      end
      12'b100101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2393;
      end
      12'b100101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2394;
      end
      12'b100101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2395;
      end
      12'b100101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2396;
      end
      12'b100101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2397;
      end
      12'b100101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2398;
      end
      12'b100101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2399;
      end
      12'b100101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2400;
      end
      12'b100101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2401;
      end
      12'b100101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2402;
      end
      12'b100101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2403;
      end
      12'b100101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2404;
      end
      12'b100101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2405;
      end
      12'b100101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2406;
      end
      12'b100101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2407;
      end
      12'b100101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2408;
      end
      12'b100101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2409;
      end
      12'b100101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2410;
      end
      12'b100101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2411;
      end
      12'b100101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2412;
      end
      12'b100101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2413;
      end
      12'b100101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2414;
      end
      12'b100101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2415;
      end
      12'b100101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2416;
      end
      12'b100101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2417;
      end
      12'b100101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2418;
      end
      12'b100101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2419;
      end
      12'b100101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2420;
      end
      12'b100101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2421;
      end
      12'b100101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2422;
      end
      12'b100101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2423;
      end
      12'b100101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2424;
      end
      12'b100101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2425;
      end
      12'b100101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2426;
      end
      12'b100101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2427;
      end
      12'b100101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2428;
      end
      12'b100101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2429;
      end
      12'b100101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2430;
      end
      12'b100101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2431;
      end
      12'b100110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2432;
      end
      12'b100110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2433;
      end
      12'b100110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2434;
      end
      12'b100110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2435;
      end
      12'b100110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2436;
      end
      12'b100110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2437;
      end
      12'b100110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2438;
      end
      12'b100110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2439;
      end
      12'b100110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2440;
      end
      12'b100110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2441;
      end
      12'b100110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2442;
      end
      12'b100110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2443;
      end
      12'b100110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2444;
      end
      12'b100110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2445;
      end
      12'b100110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2446;
      end
      12'b100110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2447;
      end
      12'b100110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2448;
      end
      12'b100110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2449;
      end
      12'b100110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2450;
      end
      12'b100110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2451;
      end
      12'b100110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2452;
      end
      12'b100110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2453;
      end
      12'b100110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2454;
      end
      12'b100110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2455;
      end
      12'b100110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2456;
      end
      12'b100110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2457;
      end
      12'b100110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2458;
      end
      12'b100110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2459;
      end
      12'b100110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2460;
      end
      12'b100110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2461;
      end
      12'b100110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2462;
      end
      12'b100110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2463;
      end
      12'b100110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2464;
      end
      12'b100110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2465;
      end
      12'b100110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2466;
      end
      12'b100110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2467;
      end
      12'b100110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2468;
      end
      12'b100110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2469;
      end
      12'b100110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2470;
      end
      12'b100110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2471;
      end
      12'b100110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2472;
      end
      12'b100110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2473;
      end
      12'b100110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2474;
      end
      12'b100110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2475;
      end
      12'b100110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2476;
      end
      12'b100110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2477;
      end
      12'b100110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2478;
      end
      12'b100110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2479;
      end
      12'b100110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2480;
      end
      12'b100110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2481;
      end
      12'b100110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2482;
      end
      12'b100110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2483;
      end
      12'b100110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2484;
      end
      12'b100110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2485;
      end
      12'b100110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2486;
      end
      12'b100110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2487;
      end
      12'b100110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2488;
      end
      12'b100110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2489;
      end
      12'b100110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2490;
      end
      12'b100110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2491;
      end
      12'b100110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2492;
      end
      12'b100110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2493;
      end
      12'b100110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2494;
      end
      12'b100110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2495;
      end
      12'b100111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2496;
      end
      12'b100111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2497;
      end
      12'b100111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2498;
      end
      12'b100111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2499;
      end
      12'b100111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2500;
      end
      12'b100111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2501;
      end
      12'b100111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2502;
      end
      12'b100111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2503;
      end
      12'b100111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2504;
      end
      12'b100111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2505;
      end
      12'b100111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2506;
      end
      12'b100111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2507;
      end
      12'b100111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2508;
      end
      12'b100111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2509;
      end
      12'b100111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2510;
      end
      12'b100111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2511;
      end
      12'b100111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2512;
      end
      12'b100111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2513;
      end
      12'b100111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2514;
      end
      12'b100111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2515;
      end
      12'b100111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2516;
      end
      12'b100111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2517;
      end
      12'b100111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2518;
      end
      12'b100111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2519;
      end
      12'b100111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2520;
      end
      12'b100111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2521;
      end
      12'b100111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2522;
      end
      12'b100111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2523;
      end
      12'b100111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2524;
      end
      12'b100111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2525;
      end
      12'b100111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2526;
      end
      12'b100111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2527;
      end
      12'b100111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2528;
      end
      12'b100111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2529;
      end
      12'b100111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2530;
      end
      12'b100111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2531;
      end
      12'b100111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2532;
      end
      12'b100111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2533;
      end
      12'b100111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2534;
      end
      12'b100111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2535;
      end
      12'b100111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2536;
      end
      12'b100111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2537;
      end
      12'b100111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2538;
      end
      12'b100111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2539;
      end
      12'b100111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2540;
      end
      12'b100111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2541;
      end
      12'b100111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2542;
      end
      12'b100111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2543;
      end
      12'b100111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2544;
      end
      12'b100111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2545;
      end
      12'b100111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2546;
      end
      12'b100111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2547;
      end
      12'b100111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2548;
      end
      12'b100111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2549;
      end
      12'b100111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2550;
      end
      12'b100111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2551;
      end
      12'b100111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2552;
      end
      12'b100111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2553;
      end
      12'b100111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2554;
      end
      12'b100111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2555;
      end
      12'b100111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2556;
      end
      12'b100111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2557;
      end
      12'b100111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2558;
      end
      12'b100111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2559;
      end
      12'b101000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2560;
      end
      12'b101000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2561;
      end
      12'b101000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2562;
      end
      12'b101000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2563;
      end
      12'b101000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2564;
      end
      12'b101000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2565;
      end
      12'b101000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2566;
      end
      12'b101000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2567;
      end
      12'b101000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2568;
      end
      12'b101000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2569;
      end
      12'b101000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2570;
      end
      12'b101000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2571;
      end
      12'b101000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2572;
      end
      12'b101000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2573;
      end
      12'b101000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2574;
      end
      12'b101000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2575;
      end
      12'b101000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2576;
      end
      12'b101000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2577;
      end
      12'b101000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2578;
      end
      12'b101000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2579;
      end
      12'b101000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2580;
      end
      12'b101000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2581;
      end
      12'b101000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2582;
      end
      12'b101000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2583;
      end
      12'b101000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2584;
      end
      12'b101000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2585;
      end
      12'b101000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2586;
      end
      12'b101000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2587;
      end
      12'b101000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2588;
      end
      12'b101000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2589;
      end
      12'b101000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2590;
      end
      12'b101000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2591;
      end
      12'b101000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2592;
      end
      12'b101000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2593;
      end
      12'b101000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2594;
      end
      12'b101000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2595;
      end
      12'b101000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2596;
      end
      12'b101000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2597;
      end
      12'b101000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2598;
      end
      12'b101000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2599;
      end
      12'b101000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2600;
      end
      12'b101000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2601;
      end
      12'b101000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2602;
      end
      12'b101000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2603;
      end
      12'b101000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2604;
      end
      12'b101000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2605;
      end
      12'b101000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2606;
      end
      12'b101000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2607;
      end
      12'b101000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2608;
      end
      12'b101000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2609;
      end
      12'b101000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2610;
      end
      12'b101000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2611;
      end
      12'b101000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2612;
      end
      12'b101000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2613;
      end
      12'b101000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2614;
      end
      12'b101000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2615;
      end
      12'b101000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2616;
      end
      12'b101000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2617;
      end
      12'b101000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2618;
      end
      12'b101000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2619;
      end
      12'b101000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2620;
      end
      12'b101000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2621;
      end
      12'b101000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2622;
      end
      12'b101000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2623;
      end
      12'b101001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2624;
      end
      12'b101001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2625;
      end
      12'b101001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2626;
      end
      12'b101001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2627;
      end
      12'b101001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2628;
      end
      12'b101001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2629;
      end
      12'b101001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2630;
      end
      12'b101001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2631;
      end
      12'b101001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2632;
      end
      12'b101001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2633;
      end
      12'b101001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2634;
      end
      12'b101001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2635;
      end
      12'b101001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2636;
      end
      12'b101001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2637;
      end
      12'b101001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2638;
      end
      12'b101001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2639;
      end
      12'b101001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2640;
      end
      12'b101001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2641;
      end
      12'b101001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2642;
      end
      12'b101001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2643;
      end
      12'b101001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2644;
      end
      12'b101001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2645;
      end
      12'b101001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2646;
      end
      12'b101001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2647;
      end
      12'b101001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2648;
      end
      12'b101001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2649;
      end
      12'b101001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2650;
      end
      12'b101001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2651;
      end
      12'b101001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2652;
      end
      12'b101001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2653;
      end
      12'b101001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2654;
      end
      12'b101001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2655;
      end
      12'b101001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2656;
      end
      12'b101001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2657;
      end
      12'b101001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2658;
      end
      12'b101001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2659;
      end
      12'b101001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2660;
      end
      12'b101001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2661;
      end
      12'b101001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2662;
      end
      12'b101001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2663;
      end
      12'b101001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2664;
      end
      12'b101001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2665;
      end
      12'b101001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2666;
      end
      12'b101001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2667;
      end
      12'b101001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2668;
      end
      12'b101001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2669;
      end
      12'b101001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2670;
      end
      12'b101001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2671;
      end
      12'b101001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2672;
      end
      12'b101001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2673;
      end
      12'b101001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2674;
      end
      12'b101001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2675;
      end
      12'b101001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2676;
      end
      12'b101001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2677;
      end
      12'b101001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2678;
      end
      12'b101001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2679;
      end
      12'b101001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2680;
      end
      12'b101001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2681;
      end
      12'b101001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2682;
      end
      12'b101001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2683;
      end
      12'b101001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2684;
      end
      12'b101001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2685;
      end
      12'b101001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2686;
      end
      12'b101001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2687;
      end
      12'b101010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2688;
      end
      12'b101010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2689;
      end
      12'b101010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2690;
      end
      12'b101010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2691;
      end
      12'b101010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2692;
      end
      12'b101010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2693;
      end
      12'b101010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2694;
      end
      12'b101010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2695;
      end
      12'b101010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2696;
      end
      12'b101010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2697;
      end
      12'b101010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2698;
      end
      12'b101010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2699;
      end
      12'b101010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2700;
      end
      12'b101010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2701;
      end
      12'b101010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2702;
      end
      12'b101010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2703;
      end
      12'b101010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2704;
      end
      12'b101010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2705;
      end
      12'b101010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2706;
      end
      12'b101010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2707;
      end
      12'b101010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2708;
      end
      12'b101010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2709;
      end
      12'b101010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2710;
      end
      12'b101010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2711;
      end
      12'b101010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2712;
      end
      12'b101010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2713;
      end
      12'b101010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2714;
      end
      12'b101010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2715;
      end
      12'b101010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2716;
      end
      12'b101010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2717;
      end
      12'b101010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2718;
      end
      12'b101010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2719;
      end
      12'b101010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2720;
      end
      12'b101010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2721;
      end
      12'b101010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2722;
      end
      12'b101010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2723;
      end
      12'b101010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2724;
      end
      12'b101010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2725;
      end
      12'b101010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2726;
      end
      12'b101010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2727;
      end
      12'b101010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2728;
      end
      12'b101010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2729;
      end
      12'b101010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2730;
      end
      12'b101010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2731;
      end
      12'b101010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2732;
      end
      12'b101010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2733;
      end
      12'b101010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2734;
      end
      12'b101010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2735;
      end
      12'b101010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2736;
      end
      12'b101010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2737;
      end
      12'b101010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2738;
      end
      12'b101010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2739;
      end
      12'b101010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2740;
      end
      12'b101010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2741;
      end
      12'b101010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2742;
      end
      12'b101010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2743;
      end
      12'b101010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2744;
      end
      12'b101010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2745;
      end
      12'b101010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2746;
      end
      12'b101010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2747;
      end
      12'b101010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2748;
      end
      12'b101010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2749;
      end
      12'b101010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2750;
      end
      12'b101010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2751;
      end
      12'b101011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2752;
      end
      12'b101011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2753;
      end
      12'b101011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2754;
      end
      12'b101011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2755;
      end
      12'b101011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2756;
      end
      12'b101011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2757;
      end
      12'b101011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2758;
      end
      12'b101011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2759;
      end
      12'b101011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2760;
      end
      12'b101011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2761;
      end
      12'b101011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2762;
      end
      12'b101011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2763;
      end
      12'b101011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2764;
      end
      12'b101011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2765;
      end
      12'b101011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2766;
      end
      12'b101011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2767;
      end
      12'b101011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2768;
      end
      12'b101011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2769;
      end
      12'b101011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2770;
      end
      12'b101011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2771;
      end
      12'b101011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2772;
      end
      12'b101011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2773;
      end
      12'b101011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2774;
      end
      12'b101011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2775;
      end
      12'b101011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2776;
      end
      12'b101011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2777;
      end
      12'b101011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2778;
      end
      12'b101011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2779;
      end
      12'b101011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2780;
      end
      12'b101011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2781;
      end
      12'b101011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2782;
      end
      12'b101011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2783;
      end
      12'b101011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2784;
      end
      12'b101011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2785;
      end
      12'b101011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2786;
      end
      12'b101011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2787;
      end
      12'b101011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2788;
      end
      12'b101011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2789;
      end
      12'b101011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2790;
      end
      12'b101011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2791;
      end
      12'b101011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2792;
      end
      12'b101011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2793;
      end
      12'b101011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2794;
      end
      12'b101011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2795;
      end
      12'b101011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2796;
      end
      12'b101011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2797;
      end
      12'b101011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2798;
      end
      12'b101011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2799;
      end
      12'b101011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2800;
      end
      12'b101011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2801;
      end
      12'b101011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2802;
      end
      12'b101011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2803;
      end
      12'b101011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2804;
      end
      12'b101011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2805;
      end
      12'b101011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2806;
      end
      12'b101011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2807;
      end
      12'b101011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2808;
      end
      12'b101011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2809;
      end
      12'b101011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2810;
      end
      12'b101011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2811;
      end
      12'b101011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2812;
      end
      12'b101011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2813;
      end
      12'b101011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2814;
      end
      12'b101011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2815;
      end
      12'b101100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2816;
      end
      12'b101100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2817;
      end
      12'b101100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2818;
      end
      12'b101100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2819;
      end
      12'b101100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2820;
      end
      12'b101100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2821;
      end
      12'b101100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2822;
      end
      12'b101100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2823;
      end
      12'b101100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2824;
      end
      12'b101100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2825;
      end
      12'b101100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2826;
      end
      12'b101100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2827;
      end
      12'b101100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2828;
      end
      12'b101100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2829;
      end
      12'b101100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2830;
      end
      12'b101100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2831;
      end
      12'b101100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2832;
      end
      12'b101100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2833;
      end
      12'b101100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2834;
      end
      12'b101100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2835;
      end
      12'b101100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2836;
      end
      12'b101100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2837;
      end
      12'b101100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2838;
      end
      12'b101100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2839;
      end
      12'b101100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2840;
      end
      12'b101100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2841;
      end
      12'b101100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2842;
      end
      12'b101100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2843;
      end
      12'b101100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2844;
      end
      12'b101100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2845;
      end
      12'b101100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2846;
      end
      12'b101100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2847;
      end
      12'b101100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2848;
      end
      12'b101100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2849;
      end
      12'b101100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2850;
      end
      12'b101100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2851;
      end
      12'b101100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2852;
      end
      12'b101100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2853;
      end
      12'b101100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2854;
      end
      12'b101100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2855;
      end
      12'b101100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2856;
      end
      12'b101100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2857;
      end
      12'b101100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2858;
      end
      12'b101100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2859;
      end
      12'b101100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2860;
      end
      12'b101100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2861;
      end
      12'b101100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2862;
      end
      12'b101100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2863;
      end
      12'b101100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2864;
      end
      12'b101100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2865;
      end
      12'b101100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2866;
      end
      12'b101100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2867;
      end
      12'b101100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2868;
      end
      12'b101100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2869;
      end
      12'b101100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2870;
      end
      12'b101100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2871;
      end
      12'b101100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2872;
      end
      12'b101100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2873;
      end
      12'b101100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2874;
      end
      12'b101100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2875;
      end
      12'b101100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2876;
      end
      12'b101100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2877;
      end
      12'b101100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2878;
      end
      12'b101100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2879;
      end
      12'b101101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2880;
      end
      12'b101101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2881;
      end
      12'b101101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2882;
      end
      12'b101101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2883;
      end
      12'b101101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2884;
      end
      12'b101101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2885;
      end
      12'b101101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2886;
      end
      12'b101101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2887;
      end
      12'b101101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2888;
      end
      12'b101101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2889;
      end
      12'b101101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2890;
      end
      12'b101101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2891;
      end
      12'b101101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2892;
      end
      12'b101101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2893;
      end
      12'b101101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2894;
      end
      12'b101101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2895;
      end
      12'b101101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2896;
      end
      12'b101101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2897;
      end
      12'b101101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2898;
      end
      12'b101101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2899;
      end
      12'b101101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2900;
      end
      12'b101101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2901;
      end
      12'b101101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2902;
      end
      12'b101101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2903;
      end
      12'b101101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2904;
      end
      12'b101101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2905;
      end
      12'b101101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2906;
      end
      12'b101101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2907;
      end
      12'b101101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2908;
      end
      12'b101101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2909;
      end
      12'b101101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2910;
      end
      12'b101101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2911;
      end
      12'b101101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2912;
      end
      12'b101101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2913;
      end
      12'b101101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2914;
      end
      12'b101101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2915;
      end
      12'b101101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2916;
      end
      12'b101101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2917;
      end
      12'b101101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2918;
      end
      12'b101101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2919;
      end
      12'b101101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2920;
      end
      12'b101101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2921;
      end
      12'b101101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2922;
      end
      12'b101101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2923;
      end
      12'b101101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2924;
      end
      12'b101101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2925;
      end
      12'b101101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2926;
      end
      12'b101101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2927;
      end
      12'b101101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2928;
      end
      12'b101101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2929;
      end
      12'b101101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2930;
      end
      12'b101101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2931;
      end
      12'b101101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2932;
      end
      12'b101101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2933;
      end
      12'b101101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2934;
      end
      12'b101101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2935;
      end
      12'b101101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2936;
      end
      12'b101101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2937;
      end
      12'b101101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2938;
      end
      12'b101101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2939;
      end
      12'b101101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2940;
      end
      12'b101101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2941;
      end
      12'b101101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2942;
      end
      12'b101101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2943;
      end
      12'b101110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2944;
      end
      12'b101110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2945;
      end
      12'b101110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2946;
      end
      12'b101110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2947;
      end
      12'b101110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2948;
      end
      12'b101110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2949;
      end
      12'b101110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2950;
      end
      12'b101110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2951;
      end
      12'b101110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2952;
      end
      12'b101110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2953;
      end
      12'b101110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2954;
      end
      12'b101110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2955;
      end
      12'b101110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2956;
      end
      12'b101110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2957;
      end
      12'b101110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2958;
      end
      12'b101110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2959;
      end
      12'b101110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2960;
      end
      12'b101110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2961;
      end
      12'b101110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2962;
      end
      12'b101110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2963;
      end
      12'b101110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2964;
      end
      12'b101110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2965;
      end
      12'b101110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2966;
      end
      12'b101110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2967;
      end
      12'b101110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2968;
      end
      12'b101110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2969;
      end
      12'b101110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2970;
      end
      12'b101110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2971;
      end
      12'b101110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2972;
      end
      12'b101110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2973;
      end
      12'b101110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2974;
      end
      12'b101110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2975;
      end
      12'b101110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2976;
      end
      12'b101110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2977;
      end
      12'b101110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2978;
      end
      12'b101110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2979;
      end
      12'b101110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2980;
      end
      12'b101110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2981;
      end
      12'b101110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2982;
      end
      12'b101110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2983;
      end
      12'b101110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2984;
      end
      12'b101110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2985;
      end
      12'b101110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2986;
      end
      12'b101110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2987;
      end
      12'b101110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2988;
      end
      12'b101110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2989;
      end
      12'b101110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2990;
      end
      12'b101110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2991;
      end
      12'b101110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_2992;
      end
      12'b101110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_2993;
      end
      12'b101110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_2994;
      end
      12'b101110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_2995;
      end
      12'b101110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_2996;
      end
      12'b101110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_2997;
      end
      12'b101110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_2998;
      end
      12'b101110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_2999;
      end
      12'b101110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3000;
      end
      12'b101110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3001;
      end
      12'b101110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3002;
      end
      12'b101110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3003;
      end
      12'b101110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3004;
      end
      12'b101110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3005;
      end
      12'b101110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3006;
      end
      12'b101110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3007;
      end
      12'b101111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3008;
      end
      12'b101111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3009;
      end
      12'b101111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3010;
      end
      12'b101111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3011;
      end
      12'b101111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3012;
      end
      12'b101111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3013;
      end
      12'b101111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3014;
      end
      12'b101111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3015;
      end
      12'b101111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3016;
      end
      12'b101111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3017;
      end
      12'b101111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3018;
      end
      12'b101111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3019;
      end
      12'b101111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3020;
      end
      12'b101111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3021;
      end
      12'b101111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3022;
      end
      12'b101111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3023;
      end
      12'b101111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3024;
      end
      12'b101111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3025;
      end
      12'b101111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3026;
      end
      12'b101111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3027;
      end
      12'b101111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3028;
      end
      12'b101111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3029;
      end
      12'b101111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3030;
      end
      12'b101111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3031;
      end
      12'b101111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3032;
      end
      12'b101111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3033;
      end
      12'b101111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3034;
      end
      12'b101111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3035;
      end
      12'b101111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3036;
      end
      12'b101111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3037;
      end
      12'b101111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3038;
      end
      12'b101111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3039;
      end
      12'b101111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3040;
      end
      12'b101111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3041;
      end
      12'b101111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3042;
      end
      12'b101111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3043;
      end
      12'b101111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3044;
      end
      12'b101111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3045;
      end
      12'b101111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3046;
      end
      12'b101111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3047;
      end
      12'b101111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3048;
      end
      12'b101111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3049;
      end
      12'b101111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3050;
      end
      12'b101111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3051;
      end
      12'b101111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3052;
      end
      12'b101111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3053;
      end
      12'b101111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3054;
      end
      12'b101111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3055;
      end
      12'b101111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3056;
      end
      12'b101111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3057;
      end
      12'b101111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3058;
      end
      12'b101111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3059;
      end
      12'b101111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3060;
      end
      12'b101111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3061;
      end
      12'b101111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3062;
      end
      12'b101111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3063;
      end
      12'b101111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3064;
      end
      12'b101111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3065;
      end
      12'b101111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3066;
      end
      12'b101111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3067;
      end
      12'b101111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3068;
      end
      12'b101111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3069;
      end
      12'b101111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3070;
      end
      12'b101111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3071;
      end
      12'b110000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3072;
      end
      12'b110000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3073;
      end
      12'b110000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3074;
      end
      12'b110000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3075;
      end
      12'b110000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3076;
      end
      12'b110000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3077;
      end
      12'b110000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3078;
      end
      12'b110000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3079;
      end
      12'b110000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3080;
      end
      12'b110000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3081;
      end
      12'b110000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3082;
      end
      12'b110000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3083;
      end
      12'b110000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3084;
      end
      12'b110000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3085;
      end
      12'b110000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3086;
      end
      12'b110000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3087;
      end
      12'b110000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3088;
      end
      12'b110000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3089;
      end
      12'b110000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3090;
      end
      12'b110000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3091;
      end
      12'b110000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3092;
      end
      12'b110000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3093;
      end
      12'b110000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3094;
      end
      12'b110000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3095;
      end
      12'b110000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3096;
      end
      12'b110000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3097;
      end
      12'b110000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3098;
      end
      12'b110000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3099;
      end
      12'b110000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3100;
      end
      12'b110000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3101;
      end
      12'b110000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3102;
      end
      12'b110000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3103;
      end
      12'b110000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3104;
      end
      12'b110000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3105;
      end
      12'b110000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3106;
      end
      12'b110000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3107;
      end
      12'b110000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3108;
      end
      12'b110000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3109;
      end
      12'b110000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3110;
      end
      12'b110000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3111;
      end
      12'b110000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3112;
      end
      12'b110000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3113;
      end
      12'b110000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3114;
      end
      12'b110000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3115;
      end
      12'b110000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3116;
      end
      12'b110000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3117;
      end
      12'b110000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3118;
      end
      12'b110000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3119;
      end
      12'b110000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3120;
      end
      12'b110000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3121;
      end
      12'b110000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3122;
      end
      12'b110000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3123;
      end
      12'b110000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3124;
      end
      12'b110000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3125;
      end
      12'b110000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3126;
      end
      12'b110000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3127;
      end
      12'b110000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3128;
      end
      12'b110000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3129;
      end
      12'b110000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3130;
      end
      12'b110000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3131;
      end
      12'b110000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3132;
      end
      12'b110000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3133;
      end
      12'b110000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3134;
      end
      12'b110000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3135;
      end
      12'b110001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3136;
      end
      12'b110001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3137;
      end
      12'b110001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3138;
      end
      12'b110001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3139;
      end
      12'b110001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3140;
      end
      12'b110001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3141;
      end
      12'b110001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3142;
      end
      12'b110001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3143;
      end
      12'b110001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3144;
      end
      12'b110001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3145;
      end
      12'b110001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3146;
      end
      12'b110001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3147;
      end
      12'b110001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3148;
      end
      12'b110001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3149;
      end
      12'b110001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3150;
      end
      12'b110001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3151;
      end
      12'b110001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3152;
      end
      12'b110001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3153;
      end
      12'b110001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3154;
      end
      12'b110001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3155;
      end
      12'b110001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3156;
      end
      12'b110001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3157;
      end
      12'b110001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3158;
      end
      12'b110001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3159;
      end
      12'b110001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3160;
      end
      12'b110001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3161;
      end
      12'b110001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3162;
      end
      12'b110001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3163;
      end
      12'b110001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3164;
      end
      12'b110001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3165;
      end
      12'b110001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3166;
      end
      12'b110001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3167;
      end
      12'b110001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3168;
      end
      12'b110001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3169;
      end
      12'b110001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3170;
      end
      12'b110001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3171;
      end
      12'b110001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3172;
      end
      12'b110001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3173;
      end
      12'b110001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3174;
      end
      12'b110001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3175;
      end
      12'b110001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3176;
      end
      12'b110001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3177;
      end
      12'b110001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3178;
      end
      12'b110001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3179;
      end
      12'b110001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3180;
      end
      12'b110001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3181;
      end
      12'b110001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3182;
      end
      12'b110001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3183;
      end
      12'b110001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3184;
      end
      12'b110001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3185;
      end
      12'b110001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3186;
      end
      12'b110001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3187;
      end
      12'b110001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3188;
      end
      12'b110001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3189;
      end
      12'b110001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3190;
      end
      12'b110001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3191;
      end
      12'b110001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3192;
      end
      12'b110001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3193;
      end
      12'b110001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3194;
      end
      12'b110001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3195;
      end
      12'b110001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3196;
      end
      12'b110001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3197;
      end
      12'b110001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3198;
      end
      12'b110001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3199;
      end
      12'b110010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3200;
      end
      12'b110010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3201;
      end
      12'b110010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3202;
      end
      12'b110010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3203;
      end
      12'b110010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3204;
      end
      12'b110010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3205;
      end
      12'b110010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3206;
      end
      12'b110010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3207;
      end
      12'b110010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3208;
      end
      12'b110010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3209;
      end
      12'b110010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3210;
      end
      12'b110010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3211;
      end
      12'b110010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3212;
      end
      12'b110010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3213;
      end
      12'b110010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3214;
      end
      12'b110010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3215;
      end
      12'b110010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3216;
      end
      12'b110010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3217;
      end
      12'b110010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3218;
      end
      12'b110010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3219;
      end
      12'b110010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3220;
      end
      12'b110010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3221;
      end
      12'b110010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3222;
      end
      12'b110010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3223;
      end
      12'b110010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3224;
      end
      12'b110010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3225;
      end
      12'b110010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3226;
      end
      12'b110010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3227;
      end
      12'b110010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3228;
      end
      12'b110010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3229;
      end
      12'b110010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3230;
      end
      12'b110010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3231;
      end
      12'b110010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3232;
      end
      12'b110010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3233;
      end
      12'b110010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3234;
      end
      12'b110010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3235;
      end
      12'b110010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3236;
      end
      12'b110010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3237;
      end
      12'b110010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3238;
      end
      12'b110010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3239;
      end
      12'b110010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3240;
      end
      12'b110010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3241;
      end
      12'b110010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3242;
      end
      12'b110010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3243;
      end
      12'b110010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3244;
      end
      12'b110010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3245;
      end
      12'b110010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3246;
      end
      12'b110010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3247;
      end
      12'b110010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3248;
      end
      12'b110010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3249;
      end
      12'b110010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3250;
      end
      12'b110010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3251;
      end
      12'b110010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3252;
      end
      12'b110010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3253;
      end
      12'b110010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3254;
      end
      12'b110010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3255;
      end
      12'b110010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3256;
      end
      12'b110010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3257;
      end
      12'b110010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3258;
      end
      12'b110010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3259;
      end
      12'b110010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3260;
      end
      12'b110010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3261;
      end
      12'b110010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3262;
      end
      12'b110010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3263;
      end
      12'b110011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3264;
      end
      12'b110011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3265;
      end
      12'b110011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3266;
      end
      12'b110011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3267;
      end
      12'b110011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3268;
      end
      12'b110011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3269;
      end
      12'b110011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3270;
      end
      12'b110011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3271;
      end
      12'b110011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3272;
      end
      12'b110011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3273;
      end
      12'b110011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3274;
      end
      12'b110011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3275;
      end
      12'b110011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3276;
      end
      12'b110011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3277;
      end
      12'b110011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3278;
      end
      12'b110011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3279;
      end
      12'b110011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3280;
      end
      12'b110011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3281;
      end
      12'b110011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3282;
      end
      12'b110011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3283;
      end
      12'b110011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3284;
      end
      12'b110011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3285;
      end
      12'b110011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3286;
      end
      12'b110011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3287;
      end
      12'b110011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3288;
      end
      12'b110011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3289;
      end
      12'b110011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3290;
      end
      12'b110011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3291;
      end
      12'b110011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3292;
      end
      12'b110011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3293;
      end
      12'b110011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3294;
      end
      12'b110011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3295;
      end
      12'b110011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3296;
      end
      12'b110011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3297;
      end
      12'b110011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3298;
      end
      12'b110011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3299;
      end
      12'b110011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3300;
      end
      12'b110011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3301;
      end
      12'b110011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3302;
      end
      12'b110011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3303;
      end
      12'b110011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3304;
      end
      12'b110011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3305;
      end
      12'b110011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3306;
      end
      12'b110011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3307;
      end
      12'b110011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3308;
      end
      12'b110011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3309;
      end
      12'b110011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3310;
      end
      12'b110011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3311;
      end
      12'b110011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3312;
      end
      12'b110011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3313;
      end
      12'b110011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3314;
      end
      12'b110011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3315;
      end
      12'b110011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3316;
      end
      12'b110011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3317;
      end
      12'b110011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3318;
      end
      12'b110011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3319;
      end
      12'b110011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3320;
      end
      12'b110011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3321;
      end
      12'b110011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3322;
      end
      12'b110011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3323;
      end
      12'b110011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3324;
      end
      12'b110011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3325;
      end
      12'b110011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3326;
      end
      12'b110011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3327;
      end
      12'b110100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3328;
      end
      12'b110100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3329;
      end
      12'b110100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3330;
      end
      12'b110100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3331;
      end
      12'b110100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3332;
      end
      12'b110100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3333;
      end
      12'b110100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3334;
      end
      12'b110100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3335;
      end
      12'b110100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3336;
      end
      12'b110100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3337;
      end
      12'b110100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3338;
      end
      12'b110100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3339;
      end
      12'b110100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3340;
      end
      12'b110100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3341;
      end
      12'b110100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3342;
      end
      12'b110100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3343;
      end
      12'b110100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3344;
      end
      12'b110100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3345;
      end
      12'b110100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3346;
      end
      12'b110100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3347;
      end
      12'b110100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3348;
      end
      12'b110100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3349;
      end
      12'b110100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3350;
      end
      12'b110100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3351;
      end
      12'b110100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3352;
      end
      12'b110100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3353;
      end
      12'b110100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3354;
      end
      12'b110100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3355;
      end
      12'b110100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3356;
      end
      12'b110100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3357;
      end
      12'b110100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3358;
      end
      12'b110100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3359;
      end
      12'b110100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3360;
      end
      12'b110100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3361;
      end
      12'b110100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3362;
      end
      12'b110100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3363;
      end
      12'b110100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3364;
      end
      12'b110100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3365;
      end
      12'b110100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3366;
      end
      12'b110100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3367;
      end
      12'b110100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3368;
      end
      12'b110100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3369;
      end
      12'b110100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3370;
      end
      12'b110100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3371;
      end
      12'b110100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3372;
      end
      12'b110100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3373;
      end
      12'b110100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3374;
      end
      12'b110100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3375;
      end
      12'b110100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3376;
      end
      12'b110100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3377;
      end
      12'b110100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3378;
      end
      12'b110100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3379;
      end
      12'b110100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3380;
      end
      12'b110100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3381;
      end
      12'b110100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3382;
      end
      12'b110100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3383;
      end
      12'b110100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3384;
      end
      12'b110100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3385;
      end
      12'b110100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3386;
      end
      12'b110100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3387;
      end
      12'b110100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3388;
      end
      12'b110100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3389;
      end
      12'b110100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3390;
      end
      12'b110100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3391;
      end
      12'b110101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3392;
      end
      12'b110101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3393;
      end
      12'b110101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3394;
      end
      12'b110101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3395;
      end
      12'b110101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3396;
      end
      12'b110101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3397;
      end
      12'b110101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3398;
      end
      12'b110101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3399;
      end
      12'b110101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3400;
      end
      12'b110101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3401;
      end
      12'b110101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3402;
      end
      12'b110101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3403;
      end
      12'b110101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3404;
      end
      12'b110101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3405;
      end
      12'b110101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3406;
      end
      12'b110101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3407;
      end
      12'b110101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3408;
      end
      12'b110101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3409;
      end
      12'b110101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3410;
      end
      12'b110101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3411;
      end
      12'b110101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3412;
      end
      12'b110101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3413;
      end
      12'b110101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3414;
      end
      12'b110101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3415;
      end
      12'b110101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3416;
      end
      12'b110101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3417;
      end
      12'b110101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3418;
      end
      12'b110101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3419;
      end
      12'b110101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3420;
      end
      12'b110101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3421;
      end
      12'b110101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3422;
      end
      12'b110101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3423;
      end
      12'b110101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3424;
      end
      12'b110101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3425;
      end
      12'b110101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3426;
      end
      12'b110101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3427;
      end
      12'b110101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3428;
      end
      12'b110101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3429;
      end
      12'b110101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3430;
      end
      12'b110101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3431;
      end
      12'b110101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3432;
      end
      12'b110101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3433;
      end
      12'b110101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3434;
      end
      12'b110101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3435;
      end
      12'b110101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3436;
      end
      12'b110101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3437;
      end
      12'b110101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3438;
      end
      12'b110101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3439;
      end
      12'b110101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3440;
      end
      12'b110101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3441;
      end
      12'b110101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3442;
      end
      12'b110101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3443;
      end
      12'b110101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3444;
      end
      12'b110101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3445;
      end
      12'b110101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3446;
      end
      12'b110101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3447;
      end
      12'b110101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3448;
      end
      12'b110101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3449;
      end
      12'b110101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3450;
      end
      12'b110101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3451;
      end
      12'b110101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3452;
      end
      12'b110101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3453;
      end
      12'b110101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3454;
      end
      12'b110101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3455;
      end
      12'b110110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3456;
      end
      12'b110110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3457;
      end
      12'b110110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3458;
      end
      12'b110110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3459;
      end
      12'b110110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3460;
      end
      12'b110110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3461;
      end
      12'b110110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3462;
      end
      12'b110110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3463;
      end
      12'b110110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3464;
      end
      12'b110110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3465;
      end
      12'b110110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3466;
      end
      12'b110110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3467;
      end
      12'b110110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3468;
      end
      12'b110110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3469;
      end
      12'b110110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3470;
      end
      12'b110110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3471;
      end
      12'b110110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3472;
      end
      12'b110110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3473;
      end
      12'b110110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3474;
      end
      12'b110110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3475;
      end
      12'b110110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3476;
      end
      12'b110110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3477;
      end
      12'b110110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3478;
      end
      12'b110110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3479;
      end
      12'b110110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3480;
      end
      12'b110110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3481;
      end
      12'b110110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3482;
      end
      12'b110110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3483;
      end
      12'b110110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3484;
      end
      12'b110110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3485;
      end
      12'b110110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3486;
      end
      12'b110110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3487;
      end
      12'b110110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3488;
      end
      12'b110110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3489;
      end
      12'b110110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3490;
      end
      12'b110110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3491;
      end
      12'b110110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3492;
      end
      12'b110110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3493;
      end
      12'b110110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3494;
      end
      12'b110110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3495;
      end
      12'b110110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3496;
      end
      12'b110110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3497;
      end
      12'b110110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3498;
      end
      12'b110110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3499;
      end
      12'b110110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3500;
      end
      12'b110110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3501;
      end
      12'b110110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3502;
      end
      12'b110110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3503;
      end
      12'b110110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3504;
      end
      12'b110110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3505;
      end
      12'b110110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3506;
      end
      12'b110110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3507;
      end
      12'b110110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3508;
      end
      12'b110110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3509;
      end
      12'b110110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3510;
      end
      12'b110110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3511;
      end
      12'b110110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3512;
      end
      12'b110110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3513;
      end
      12'b110110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3514;
      end
      12'b110110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3515;
      end
      12'b110110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3516;
      end
      12'b110110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3517;
      end
      12'b110110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3518;
      end
      12'b110110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3519;
      end
      12'b110111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3520;
      end
      12'b110111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3521;
      end
      12'b110111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3522;
      end
      12'b110111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3523;
      end
      12'b110111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3524;
      end
      12'b110111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3525;
      end
      12'b110111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3526;
      end
      12'b110111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3527;
      end
      12'b110111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3528;
      end
      12'b110111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3529;
      end
      12'b110111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3530;
      end
      12'b110111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3531;
      end
      12'b110111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3532;
      end
      12'b110111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3533;
      end
      12'b110111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3534;
      end
      12'b110111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3535;
      end
      12'b110111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3536;
      end
      12'b110111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3537;
      end
      12'b110111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3538;
      end
      12'b110111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3539;
      end
      12'b110111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3540;
      end
      12'b110111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3541;
      end
      12'b110111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3542;
      end
      12'b110111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3543;
      end
      12'b110111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3544;
      end
      12'b110111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3545;
      end
      12'b110111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3546;
      end
      12'b110111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3547;
      end
      12'b110111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3548;
      end
      12'b110111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3549;
      end
      12'b110111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3550;
      end
      12'b110111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3551;
      end
      12'b110111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3552;
      end
      12'b110111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3553;
      end
      12'b110111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3554;
      end
      12'b110111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3555;
      end
      12'b110111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3556;
      end
      12'b110111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3557;
      end
      12'b110111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3558;
      end
      12'b110111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3559;
      end
      12'b110111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3560;
      end
      12'b110111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3561;
      end
      12'b110111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3562;
      end
      12'b110111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3563;
      end
      12'b110111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3564;
      end
      12'b110111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3565;
      end
      12'b110111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3566;
      end
      12'b110111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3567;
      end
      12'b110111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3568;
      end
      12'b110111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3569;
      end
      12'b110111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3570;
      end
      12'b110111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3571;
      end
      12'b110111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3572;
      end
      12'b110111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3573;
      end
      12'b110111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3574;
      end
      12'b110111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3575;
      end
      12'b110111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3576;
      end
      12'b110111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3577;
      end
      12'b110111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3578;
      end
      12'b110111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3579;
      end
      12'b110111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3580;
      end
      12'b110111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3581;
      end
      12'b110111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3582;
      end
      12'b110111111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3583;
      end
      12'b111000000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3584;
      end
      12'b111000000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3585;
      end
      12'b111000000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3586;
      end
      12'b111000000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3587;
      end
      12'b111000000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3588;
      end
      12'b111000000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3589;
      end
      12'b111000000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3590;
      end
      12'b111000000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3591;
      end
      12'b111000001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3592;
      end
      12'b111000001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3593;
      end
      12'b111000001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3594;
      end
      12'b111000001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3595;
      end
      12'b111000001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3596;
      end
      12'b111000001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3597;
      end
      12'b111000001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3598;
      end
      12'b111000001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3599;
      end
      12'b111000010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3600;
      end
      12'b111000010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3601;
      end
      12'b111000010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3602;
      end
      12'b111000010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3603;
      end
      12'b111000010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3604;
      end
      12'b111000010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3605;
      end
      12'b111000010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3606;
      end
      12'b111000010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3607;
      end
      12'b111000011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3608;
      end
      12'b111000011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3609;
      end
      12'b111000011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3610;
      end
      12'b111000011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3611;
      end
      12'b111000011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3612;
      end
      12'b111000011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3613;
      end
      12'b111000011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3614;
      end
      12'b111000011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3615;
      end
      12'b111000100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3616;
      end
      12'b111000100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3617;
      end
      12'b111000100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3618;
      end
      12'b111000100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3619;
      end
      12'b111000100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3620;
      end
      12'b111000100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3621;
      end
      12'b111000100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3622;
      end
      12'b111000100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3623;
      end
      12'b111000101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3624;
      end
      12'b111000101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3625;
      end
      12'b111000101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3626;
      end
      12'b111000101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3627;
      end
      12'b111000101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3628;
      end
      12'b111000101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3629;
      end
      12'b111000101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3630;
      end
      12'b111000101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3631;
      end
      12'b111000110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3632;
      end
      12'b111000110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3633;
      end
      12'b111000110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3634;
      end
      12'b111000110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3635;
      end
      12'b111000110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3636;
      end
      12'b111000110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3637;
      end
      12'b111000110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3638;
      end
      12'b111000110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3639;
      end
      12'b111000111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3640;
      end
      12'b111000111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3641;
      end
      12'b111000111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3642;
      end
      12'b111000111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3643;
      end
      12'b111000111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3644;
      end
      12'b111000111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3645;
      end
      12'b111000111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3646;
      end
      12'b111000111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3647;
      end
      12'b111001000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3648;
      end
      12'b111001000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3649;
      end
      12'b111001000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3650;
      end
      12'b111001000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3651;
      end
      12'b111001000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3652;
      end
      12'b111001000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3653;
      end
      12'b111001000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3654;
      end
      12'b111001000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3655;
      end
      12'b111001001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3656;
      end
      12'b111001001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3657;
      end
      12'b111001001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3658;
      end
      12'b111001001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3659;
      end
      12'b111001001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3660;
      end
      12'b111001001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3661;
      end
      12'b111001001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3662;
      end
      12'b111001001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3663;
      end
      12'b111001010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3664;
      end
      12'b111001010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3665;
      end
      12'b111001010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3666;
      end
      12'b111001010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3667;
      end
      12'b111001010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3668;
      end
      12'b111001010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3669;
      end
      12'b111001010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3670;
      end
      12'b111001010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3671;
      end
      12'b111001011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3672;
      end
      12'b111001011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3673;
      end
      12'b111001011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3674;
      end
      12'b111001011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3675;
      end
      12'b111001011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3676;
      end
      12'b111001011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3677;
      end
      12'b111001011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3678;
      end
      12'b111001011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3679;
      end
      12'b111001100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3680;
      end
      12'b111001100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3681;
      end
      12'b111001100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3682;
      end
      12'b111001100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3683;
      end
      12'b111001100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3684;
      end
      12'b111001100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3685;
      end
      12'b111001100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3686;
      end
      12'b111001100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3687;
      end
      12'b111001101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3688;
      end
      12'b111001101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3689;
      end
      12'b111001101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3690;
      end
      12'b111001101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3691;
      end
      12'b111001101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3692;
      end
      12'b111001101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3693;
      end
      12'b111001101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3694;
      end
      12'b111001101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3695;
      end
      12'b111001110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3696;
      end
      12'b111001110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3697;
      end
      12'b111001110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3698;
      end
      12'b111001110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3699;
      end
      12'b111001110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3700;
      end
      12'b111001110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3701;
      end
      12'b111001110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3702;
      end
      12'b111001110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3703;
      end
      12'b111001111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3704;
      end
      12'b111001111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3705;
      end
      12'b111001111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3706;
      end
      12'b111001111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3707;
      end
      12'b111001111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3708;
      end
      12'b111001111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3709;
      end
      12'b111001111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3710;
      end
      12'b111001111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3711;
      end
      12'b111010000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3712;
      end
      12'b111010000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3713;
      end
      12'b111010000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3714;
      end
      12'b111010000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3715;
      end
      12'b111010000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3716;
      end
      12'b111010000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3717;
      end
      12'b111010000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3718;
      end
      12'b111010000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3719;
      end
      12'b111010001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3720;
      end
      12'b111010001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3721;
      end
      12'b111010001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3722;
      end
      12'b111010001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3723;
      end
      12'b111010001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3724;
      end
      12'b111010001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3725;
      end
      12'b111010001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3726;
      end
      12'b111010001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3727;
      end
      12'b111010010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3728;
      end
      12'b111010010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3729;
      end
      12'b111010010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3730;
      end
      12'b111010010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3731;
      end
      12'b111010010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3732;
      end
      12'b111010010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3733;
      end
      12'b111010010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3734;
      end
      12'b111010010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3735;
      end
      12'b111010011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3736;
      end
      12'b111010011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3737;
      end
      12'b111010011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3738;
      end
      12'b111010011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3739;
      end
      12'b111010011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3740;
      end
      12'b111010011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3741;
      end
      12'b111010011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3742;
      end
      12'b111010011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3743;
      end
      12'b111010100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3744;
      end
      12'b111010100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3745;
      end
      12'b111010100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3746;
      end
      12'b111010100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3747;
      end
      12'b111010100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3748;
      end
      12'b111010100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3749;
      end
      12'b111010100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3750;
      end
      12'b111010100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3751;
      end
      12'b111010101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3752;
      end
      12'b111010101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3753;
      end
      12'b111010101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3754;
      end
      12'b111010101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3755;
      end
      12'b111010101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3756;
      end
      12'b111010101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3757;
      end
      12'b111010101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3758;
      end
      12'b111010101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3759;
      end
      12'b111010110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3760;
      end
      12'b111010110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3761;
      end
      12'b111010110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3762;
      end
      12'b111010110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3763;
      end
      12'b111010110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3764;
      end
      12'b111010110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3765;
      end
      12'b111010110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3766;
      end
      12'b111010110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3767;
      end
      12'b111010111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3768;
      end
      12'b111010111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3769;
      end
      12'b111010111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3770;
      end
      12'b111010111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3771;
      end
      12'b111010111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3772;
      end
      12'b111010111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3773;
      end
      12'b111010111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3774;
      end
      12'b111010111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3775;
      end
      12'b111011000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3776;
      end
      12'b111011000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3777;
      end
      12'b111011000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3778;
      end
      12'b111011000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3779;
      end
      12'b111011000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3780;
      end
      12'b111011000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3781;
      end
      12'b111011000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3782;
      end
      12'b111011000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3783;
      end
      12'b111011001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3784;
      end
      12'b111011001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3785;
      end
      12'b111011001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3786;
      end
      12'b111011001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3787;
      end
      12'b111011001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3788;
      end
      12'b111011001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3789;
      end
      12'b111011001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3790;
      end
      12'b111011001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3791;
      end
      12'b111011010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3792;
      end
      12'b111011010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3793;
      end
      12'b111011010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3794;
      end
      12'b111011010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3795;
      end
      12'b111011010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3796;
      end
      12'b111011010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3797;
      end
      12'b111011010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3798;
      end
      12'b111011010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3799;
      end
      12'b111011011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3800;
      end
      12'b111011011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3801;
      end
      12'b111011011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3802;
      end
      12'b111011011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3803;
      end
      12'b111011011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3804;
      end
      12'b111011011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3805;
      end
      12'b111011011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3806;
      end
      12'b111011011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3807;
      end
      12'b111011100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3808;
      end
      12'b111011100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3809;
      end
      12'b111011100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3810;
      end
      12'b111011100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3811;
      end
      12'b111011100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3812;
      end
      12'b111011100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3813;
      end
      12'b111011100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3814;
      end
      12'b111011100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3815;
      end
      12'b111011101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3816;
      end
      12'b111011101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3817;
      end
      12'b111011101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3818;
      end
      12'b111011101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3819;
      end
      12'b111011101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3820;
      end
      12'b111011101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3821;
      end
      12'b111011101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3822;
      end
      12'b111011101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3823;
      end
      12'b111011110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3824;
      end
      12'b111011110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3825;
      end
      12'b111011110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3826;
      end
      12'b111011110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3827;
      end
      12'b111011110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3828;
      end
      12'b111011110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3829;
      end
      12'b111011110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3830;
      end
      12'b111011110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3831;
      end
      12'b111011111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3832;
      end
      12'b111011111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3833;
      end
      12'b111011111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3834;
      end
      12'b111011111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3835;
      end
      12'b111011111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3836;
      end
      12'b111011111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3837;
      end
      12'b111011111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3838;
      end
      12'b111011111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3839;
      end
      12'b111100000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3840;
      end
      12'b111100000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3841;
      end
      12'b111100000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3842;
      end
      12'b111100000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3843;
      end
      12'b111100000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3844;
      end
      12'b111100000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3845;
      end
      12'b111100000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3846;
      end
      12'b111100000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3847;
      end
      12'b111100001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3848;
      end
      12'b111100001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3849;
      end
      12'b111100001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3850;
      end
      12'b111100001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3851;
      end
      12'b111100001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3852;
      end
      12'b111100001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3853;
      end
      12'b111100001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3854;
      end
      12'b111100001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3855;
      end
      12'b111100010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3856;
      end
      12'b111100010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3857;
      end
      12'b111100010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3858;
      end
      12'b111100010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3859;
      end
      12'b111100010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3860;
      end
      12'b111100010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3861;
      end
      12'b111100010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3862;
      end
      12'b111100010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3863;
      end
      12'b111100011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3864;
      end
      12'b111100011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3865;
      end
      12'b111100011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3866;
      end
      12'b111100011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3867;
      end
      12'b111100011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3868;
      end
      12'b111100011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3869;
      end
      12'b111100011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3870;
      end
      12'b111100011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3871;
      end
      12'b111100100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3872;
      end
      12'b111100100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3873;
      end
      12'b111100100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3874;
      end
      12'b111100100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3875;
      end
      12'b111100100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3876;
      end
      12'b111100100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3877;
      end
      12'b111100100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3878;
      end
      12'b111100100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3879;
      end
      12'b111100101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3880;
      end
      12'b111100101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3881;
      end
      12'b111100101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3882;
      end
      12'b111100101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3883;
      end
      12'b111100101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3884;
      end
      12'b111100101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3885;
      end
      12'b111100101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3886;
      end
      12'b111100101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3887;
      end
      12'b111100110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3888;
      end
      12'b111100110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3889;
      end
      12'b111100110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3890;
      end
      12'b111100110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3891;
      end
      12'b111100110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3892;
      end
      12'b111100110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3893;
      end
      12'b111100110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3894;
      end
      12'b111100110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3895;
      end
      12'b111100111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3896;
      end
      12'b111100111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3897;
      end
      12'b111100111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3898;
      end
      12'b111100111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3899;
      end
      12'b111100111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3900;
      end
      12'b111100111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3901;
      end
      12'b111100111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3902;
      end
      12'b111100111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3903;
      end
      12'b111101000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3904;
      end
      12'b111101000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3905;
      end
      12'b111101000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3906;
      end
      12'b111101000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3907;
      end
      12'b111101000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3908;
      end
      12'b111101000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3909;
      end
      12'b111101000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3910;
      end
      12'b111101000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3911;
      end
      12'b111101001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3912;
      end
      12'b111101001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3913;
      end
      12'b111101001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3914;
      end
      12'b111101001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3915;
      end
      12'b111101001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3916;
      end
      12'b111101001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3917;
      end
      12'b111101001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3918;
      end
      12'b111101001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3919;
      end
      12'b111101010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3920;
      end
      12'b111101010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3921;
      end
      12'b111101010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3922;
      end
      12'b111101010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3923;
      end
      12'b111101010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3924;
      end
      12'b111101010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3925;
      end
      12'b111101010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3926;
      end
      12'b111101010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3927;
      end
      12'b111101011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3928;
      end
      12'b111101011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3929;
      end
      12'b111101011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3930;
      end
      12'b111101011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3931;
      end
      12'b111101011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3932;
      end
      12'b111101011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3933;
      end
      12'b111101011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3934;
      end
      12'b111101011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3935;
      end
      12'b111101100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3936;
      end
      12'b111101100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3937;
      end
      12'b111101100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3938;
      end
      12'b111101100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3939;
      end
      12'b111101100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3940;
      end
      12'b111101100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3941;
      end
      12'b111101100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3942;
      end
      12'b111101100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3943;
      end
      12'b111101101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3944;
      end
      12'b111101101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3945;
      end
      12'b111101101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3946;
      end
      12'b111101101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3947;
      end
      12'b111101101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3948;
      end
      12'b111101101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3949;
      end
      12'b111101101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3950;
      end
      12'b111101101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3951;
      end
      12'b111101110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3952;
      end
      12'b111101110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3953;
      end
      12'b111101110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3954;
      end
      12'b111101110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3955;
      end
      12'b111101110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3956;
      end
      12'b111101110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3957;
      end
      12'b111101110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3958;
      end
      12'b111101110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3959;
      end
      12'b111101111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3960;
      end
      12'b111101111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3961;
      end
      12'b111101111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3962;
      end
      12'b111101111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3963;
      end
      12'b111101111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3964;
      end
      12'b111101111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3965;
      end
      12'b111101111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3966;
      end
      12'b111101111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3967;
      end
      12'b111110000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3968;
      end
      12'b111110000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3969;
      end
      12'b111110000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3970;
      end
      12'b111110000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3971;
      end
      12'b111110000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3972;
      end
      12'b111110000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3973;
      end
      12'b111110000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3974;
      end
      12'b111110000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3975;
      end
      12'b111110001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3976;
      end
      12'b111110001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3977;
      end
      12'b111110001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3978;
      end
      12'b111110001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3979;
      end
      12'b111110001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3980;
      end
      12'b111110001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3981;
      end
      12'b111110001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3982;
      end
      12'b111110001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3983;
      end
      12'b111110010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3984;
      end
      12'b111110010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3985;
      end
      12'b111110010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3986;
      end
      12'b111110010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3987;
      end
      12'b111110010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3988;
      end
      12'b111110010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3989;
      end
      12'b111110010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3990;
      end
      12'b111110010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3991;
      end
      12'b111110011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_3992;
      end
      12'b111110011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_3993;
      end
      12'b111110011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_3994;
      end
      12'b111110011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_3995;
      end
      12'b111110011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_3996;
      end
      12'b111110011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_3997;
      end
      12'b111110011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_3998;
      end
      12'b111110011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_3999;
      end
      12'b111110100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4000;
      end
      12'b111110100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4001;
      end
      12'b111110100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4002;
      end
      12'b111110100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4003;
      end
      12'b111110100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4004;
      end
      12'b111110100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4005;
      end
      12'b111110100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4006;
      end
      12'b111110100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4007;
      end
      12'b111110101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4008;
      end
      12'b111110101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4009;
      end
      12'b111110101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4010;
      end
      12'b111110101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4011;
      end
      12'b111110101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4012;
      end
      12'b111110101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4013;
      end
      12'b111110101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4014;
      end
      12'b111110101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4015;
      end
      12'b111110110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4016;
      end
      12'b111110110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4017;
      end
      12'b111110110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4018;
      end
      12'b111110110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4019;
      end
      12'b111110110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4020;
      end
      12'b111110110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4021;
      end
      12'b111110110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4022;
      end
      12'b111110110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4023;
      end
      12'b111110111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4024;
      end
      12'b111110111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4025;
      end
      12'b111110111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4026;
      end
      12'b111110111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4027;
      end
      12'b111110111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4028;
      end
      12'b111110111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4029;
      end
      12'b111110111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4030;
      end
      12'b111110111111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4031;
      end
      12'b111111000000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4032;
      end
      12'b111111000001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4033;
      end
      12'b111111000010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4034;
      end
      12'b111111000011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4035;
      end
      12'b111111000100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4036;
      end
      12'b111111000101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4037;
      end
      12'b111111000110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4038;
      end
      12'b111111000111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4039;
      end
      12'b111111001000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4040;
      end
      12'b111111001001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4041;
      end
      12'b111111001010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4042;
      end
      12'b111111001011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4043;
      end
      12'b111111001100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4044;
      end
      12'b111111001101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4045;
      end
      12'b111111001110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4046;
      end
      12'b111111001111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4047;
      end
      12'b111111010000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4048;
      end
      12'b111111010001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4049;
      end
      12'b111111010010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4050;
      end
      12'b111111010011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4051;
      end
      12'b111111010100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4052;
      end
      12'b111111010101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4053;
      end
      12'b111111010110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4054;
      end
      12'b111111010111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4055;
      end
      12'b111111011000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4056;
      end
      12'b111111011001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4057;
      end
      12'b111111011010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4058;
      end
      12'b111111011011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4059;
      end
      12'b111111011100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4060;
      end
      12'b111111011101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4061;
      end
      12'b111111011110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4062;
      end
      12'b111111011111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4063;
      end
      12'b111111100000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4064;
      end
      12'b111111100001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4065;
      end
      12'b111111100010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4066;
      end
      12'b111111100011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4067;
      end
      12'b111111100100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4068;
      end
      12'b111111100101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4069;
      end
      12'b111111100110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4070;
      end
      12'b111111100111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4071;
      end
      12'b111111101000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4072;
      end
      12'b111111101001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4073;
      end
      12'b111111101010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4074;
      end
      12'b111111101011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4075;
      end
      12'b111111101100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4076;
      end
      12'b111111101101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4077;
      end
      12'b111111101110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4078;
      end
      12'b111111101111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4079;
      end
      12'b111111110000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4080;
      end
      12'b111111110001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4081;
      end
      12'b111111110010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4082;
      end
      12'b111111110011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4083;
      end
      12'b111111110100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4084;
      end
      12'b111111110101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4085;
      end
      12'b111111110110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4086;
      end
      12'b111111110111 : begin
        _zz__zz_regVec_0_1_1 = regVec_4087;
      end
      12'b111111111000 : begin
        _zz__zz_regVec_0_1_1 = regVec_4088;
      end
      12'b111111111001 : begin
        _zz__zz_regVec_0_1_1 = regVec_4089;
      end
      12'b111111111010 : begin
        _zz__zz_regVec_0_1_1 = regVec_4090;
      end
      12'b111111111011 : begin
        _zz__zz_regVec_0_1_1 = regVec_4091;
      end
      12'b111111111100 : begin
        _zz__zz_regVec_0_1_1 = regVec_4092;
      end
      12'b111111111101 : begin
        _zz__zz_regVec_0_1_1 = regVec_4093;
      end
      12'b111111111110 : begin
        _zz__zz_regVec_0_1_1 = regVec_4094;
      end
      default : begin
        _zz__zz_regVec_0_1_1 = regVec_4095;
      end
    endcase
  end

  always @(*) begin
    case(Axi4Incr_wrapCase)
      2'b00 : begin
        _zz_Axi4Incr_result = {Axi4Incr_base[11 : 1],Axi4Incr_baseIncr[0 : 0]};
      end
      2'b01 : begin
        _zz_Axi4Incr_result = {Axi4Incr_base[11 : 2],Axi4Incr_baseIncr[1 : 0]};
      end
      2'b10 : begin
        _zz_Axi4Incr_result = {Axi4Incr_base[11 : 3],Axi4Incr_baseIncr[2 : 0]};
      end
      default : begin
        _zz_Axi4Incr_result = {Axi4Incr_base[11 : 4],Axi4Incr_baseIncr[3 : 0]};
      end
    endcase
  end

  always @(*) begin
    case(_zz_axiSignal_r_payload_data_1)
      12'b000000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_0;
      end
      12'b000000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1;
      end
      12'b000000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2;
      end
      12'b000000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3;
      end
      12'b000000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_4;
      end
      12'b000000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_5;
      end
      12'b000000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_6;
      end
      12'b000000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_7;
      end
      12'b000000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_8;
      end
      12'b000000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_9;
      end
      12'b000000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_10;
      end
      12'b000000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_11;
      end
      12'b000000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_12;
      end
      12'b000000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_13;
      end
      12'b000000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_14;
      end
      12'b000000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_15;
      end
      12'b000000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_16;
      end
      12'b000000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_17;
      end
      12'b000000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_18;
      end
      12'b000000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_19;
      end
      12'b000000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_20;
      end
      12'b000000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_21;
      end
      12'b000000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_22;
      end
      12'b000000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_23;
      end
      12'b000000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_24;
      end
      12'b000000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_25;
      end
      12'b000000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_26;
      end
      12'b000000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_27;
      end
      12'b000000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_28;
      end
      12'b000000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_29;
      end
      12'b000000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_30;
      end
      12'b000000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_31;
      end
      12'b000000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_32;
      end
      12'b000000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_33;
      end
      12'b000000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_34;
      end
      12'b000000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_35;
      end
      12'b000000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_36;
      end
      12'b000000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_37;
      end
      12'b000000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_38;
      end
      12'b000000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_39;
      end
      12'b000000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_40;
      end
      12'b000000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_41;
      end
      12'b000000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_42;
      end
      12'b000000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_43;
      end
      12'b000000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_44;
      end
      12'b000000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_45;
      end
      12'b000000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_46;
      end
      12'b000000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_47;
      end
      12'b000000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_48;
      end
      12'b000000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_49;
      end
      12'b000000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_50;
      end
      12'b000000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_51;
      end
      12'b000000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_52;
      end
      12'b000000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_53;
      end
      12'b000000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_54;
      end
      12'b000000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_55;
      end
      12'b000000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_56;
      end
      12'b000000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_57;
      end
      12'b000000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_58;
      end
      12'b000000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_59;
      end
      12'b000000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_60;
      end
      12'b000000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_61;
      end
      12'b000000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_62;
      end
      12'b000000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_63;
      end
      12'b000001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_64;
      end
      12'b000001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_65;
      end
      12'b000001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_66;
      end
      12'b000001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_67;
      end
      12'b000001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_68;
      end
      12'b000001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_69;
      end
      12'b000001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_70;
      end
      12'b000001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_71;
      end
      12'b000001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_72;
      end
      12'b000001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_73;
      end
      12'b000001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_74;
      end
      12'b000001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_75;
      end
      12'b000001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_76;
      end
      12'b000001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_77;
      end
      12'b000001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_78;
      end
      12'b000001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_79;
      end
      12'b000001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_80;
      end
      12'b000001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_81;
      end
      12'b000001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_82;
      end
      12'b000001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_83;
      end
      12'b000001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_84;
      end
      12'b000001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_85;
      end
      12'b000001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_86;
      end
      12'b000001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_87;
      end
      12'b000001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_88;
      end
      12'b000001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_89;
      end
      12'b000001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_90;
      end
      12'b000001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_91;
      end
      12'b000001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_92;
      end
      12'b000001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_93;
      end
      12'b000001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_94;
      end
      12'b000001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_95;
      end
      12'b000001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_96;
      end
      12'b000001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_97;
      end
      12'b000001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_98;
      end
      12'b000001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_99;
      end
      12'b000001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_100;
      end
      12'b000001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_101;
      end
      12'b000001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_102;
      end
      12'b000001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_103;
      end
      12'b000001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_104;
      end
      12'b000001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_105;
      end
      12'b000001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_106;
      end
      12'b000001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_107;
      end
      12'b000001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_108;
      end
      12'b000001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_109;
      end
      12'b000001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_110;
      end
      12'b000001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_111;
      end
      12'b000001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_112;
      end
      12'b000001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_113;
      end
      12'b000001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_114;
      end
      12'b000001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_115;
      end
      12'b000001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_116;
      end
      12'b000001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_117;
      end
      12'b000001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_118;
      end
      12'b000001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_119;
      end
      12'b000001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_120;
      end
      12'b000001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_121;
      end
      12'b000001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_122;
      end
      12'b000001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_123;
      end
      12'b000001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_124;
      end
      12'b000001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_125;
      end
      12'b000001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_126;
      end
      12'b000001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_127;
      end
      12'b000010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_128;
      end
      12'b000010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_129;
      end
      12'b000010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_130;
      end
      12'b000010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_131;
      end
      12'b000010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_132;
      end
      12'b000010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_133;
      end
      12'b000010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_134;
      end
      12'b000010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_135;
      end
      12'b000010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_136;
      end
      12'b000010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_137;
      end
      12'b000010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_138;
      end
      12'b000010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_139;
      end
      12'b000010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_140;
      end
      12'b000010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_141;
      end
      12'b000010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_142;
      end
      12'b000010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_143;
      end
      12'b000010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_144;
      end
      12'b000010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_145;
      end
      12'b000010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_146;
      end
      12'b000010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_147;
      end
      12'b000010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_148;
      end
      12'b000010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_149;
      end
      12'b000010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_150;
      end
      12'b000010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_151;
      end
      12'b000010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_152;
      end
      12'b000010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_153;
      end
      12'b000010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_154;
      end
      12'b000010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_155;
      end
      12'b000010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_156;
      end
      12'b000010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_157;
      end
      12'b000010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_158;
      end
      12'b000010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_159;
      end
      12'b000010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_160;
      end
      12'b000010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_161;
      end
      12'b000010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_162;
      end
      12'b000010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_163;
      end
      12'b000010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_164;
      end
      12'b000010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_165;
      end
      12'b000010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_166;
      end
      12'b000010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_167;
      end
      12'b000010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_168;
      end
      12'b000010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_169;
      end
      12'b000010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_170;
      end
      12'b000010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_171;
      end
      12'b000010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_172;
      end
      12'b000010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_173;
      end
      12'b000010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_174;
      end
      12'b000010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_175;
      end
      12'b000010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_176;
      end
      12'b000010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_177;
      end
      12'b000010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_178;
      end
      12'b000010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_179;
      end
      12'b000010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_180;
      end
      12'b000010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_181;
      end
      12'b000010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_182;
      end
      12'b000010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_183;
      end
      12'b000010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_184;
      end
      12'b000010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_185;
      end
      12'b000010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_186;
      end
      12'b000010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_187;
      end
      12'b000010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_188;
      end
      12'b000010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_189;
      end
      12'b000010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_190;
      end
      12'b000010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_191;
      end
      12'b000011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_192;
      end
      12'b000011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_193;
      end
      12'b000011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_194;
      end
      12'b000011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_195;
      end
      12'b000011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_196;
      end
      12'b000011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_197;
      end
      12'b000011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_198;
      end
      12'b000011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_199;
      end
      12'b000011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_200;
      end
      12'b000011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_201;
      end
      12'b000011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_202;
      end
      12'b000011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_203;
      end
      12'b000011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_204;
      end
      12'b000011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_205;
      end
      12'b000011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_206;
      end
      12'b000011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_207;
      end
      12'b000011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_208;
      end
      12'b000011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_209;
      end
      12'b000011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_210;
      end
      12'b000011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_211;
      end
      12'b000011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_212;
      end
      12'b000011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_213;
      end
      12'b000011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_214;
      end
      12'b000011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_215;
      end
      12'b000011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_216;
      end
      12'b000011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_217;
      end
      12'b000011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_218;
      end
      12'b000011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_219;
      end
      12'b000011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_220;
      end
      12'b000011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_221;
      end
      12'b000011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_222;
      end
      12'b000011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_223;
      end
      12'b000011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_224;
      end
      12'b000011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_225;
      end
      12'b000011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_226;
      end
      12'b000011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_227;
      end
      12'b000011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_228;
      end
      12'b000011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_229;
      end
      12'b000011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_230;
      end
      12'b000011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_231;
      end
      12'b000011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_232;
      end
      12'b000011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_233;
      end
      12'b000011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_234;
      end
      12'b000011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_235;
      end
      12'b000011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_236;
      end
      12'b000011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_237;
      end
      12'b000011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_238;
      end
      12'b000011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_239;
      end
      12'b000011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_240;
      end
      12'b000011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_241;
      end
      12'b000011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_242;
      end
      12'b000011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_243;
      end
      12'b000011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_244;
      end
      12'b000011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_245;
      end
      12'b000011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_246;
      end
      12'b000011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_247;
      end
      12'b000011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_248;
      end
      12'b000011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_249;
      end
      12'b000011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_250;
      end
      12'b000011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_251;
      end
      12'b000011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_252;
      end
      12'b000011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_253;
      end
      12'b000011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_254;
      end
      12'b000011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_255;
      end
      12'b000100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_256;
      end
      12'b000100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_257;
      end
      12'b000100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_258;
      end
      12'b000100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_259;
      end
      12'b000100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_260;
      end
      12'b000100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_261;
      end
      12'b000100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_262;
      end
      12'b000100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_263;
      end
      12'b000100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_264;
      end
      12'b000100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_265;
      end
      12'b000100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_266;
      end
      12'b000100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_267;
      end
      12'b000100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_268;
      end
      12'b000100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_269;
      end
      12'b000100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_270;
      end
      12'b000100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_271;
      end
      12'b000100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_272;
      end
      12'b000100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_273;
      end
      12'b000100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_274;
      end
      12'b000100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_275;
      end
      12'b000100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_276;
      end
      12'b000100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_277;
      end
      12'b000100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_278;
      end
      12'b000100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_279;
      end
      12'b000100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_280;
      end
      12'b000100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_281;
      end
      12'b000100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_282;
      end
      12'b000100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_283;
      end
      12'b000100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_284;
      end
      12'b000100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_285;
      end
      12'b000100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_286;
      end
      12'b000100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_287;
      end
      12'b000100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_288;
      end
      12'b000100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_289;
      end
      12'b000100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_290;
      end
      12'b000100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_291;
      end
      12'b000100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_292;
      end
      12'b000100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_293;
      end
      12'b000100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_294;
      end
      12'b000100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_295;
      end
      12'b000100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_296;
      end
      12'b000100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_297;
      end
      12'b000100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_298;
      end
      12'b000100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_299;
      end
      12'b000100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_300;
      end
      12'b000100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_301;
      end
      12'b000100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_302;
      end
      12'b000100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_303;
      end
      12'b000100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_304;
      end
      12'b000100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_305;
      end
      12'b000100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_306;
      end
      12'b000100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_307;
      end
      12'b000100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_308;
      end
      12'b000100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_309;
      end
      12'b000100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_310;
      end
      12'b000100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_311;
      end
      12'b000100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_312;
      end
      12'b000100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_313;
      end
      12'b000100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_314;
      end
      12'b000100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_315;
      end
      12'b000100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_316;
      end
      12'b000100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_317;
      end
      12'b000100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_318;
      end
      12'b000100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_319;
      end
      12'b000101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_320;
      end
      12'b000101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_321;
      end
      12'b000101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_322;
      end
      12'b000101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_323;
      end
      12'b000101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_324;
      end
      12'b000101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_325;
      end
      12'b000101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_326;
      end
      12'b000101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_327;
      end
      12'b000101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_328;
      end
      12'b000101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_329;
      end
      12'b000101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_330;
      end
      12'b000101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_331;
      end
      12'b000101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_332;
      end
      12'b000101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_333;
      end
      12'b000101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_334;
      end
      12'b000101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_335;
      end
      12'b000101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_336;
      end
      12'b000101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_337;
      end
      12'b000101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_338;
      end
      12'b000101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_339;
      end
      12'b000101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_340;
      end
      12'b000101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_341;
      end
      12'b000101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_342;
      end
      12'b000101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_343;
      end
      12'b000101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_344;
      end
      12'b000101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_345;
      end
      12'b000101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_346;
      end
      12'b000101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_347;
      end
      12'b000101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_348;
      end
      12'b000101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_349;
      end
      12'b000101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_350;
      end
      12'b000101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_351;
      end
      12'b000101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_352;
      end
      12'b000101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_353;
      end
      12'b000101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_354;
      end
      12'b000101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_355;
      end
      12'b000101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_356;
      end
      12'b000101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_357;
      end
      12'b000101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_358;
      end
      12'b000101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_359;
      end
      12'b000101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_360;
      end
      12'b000101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_361;
      end
      12'b000101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_362;
      end
      12'b000101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_363;
      end
      12'b000101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_364;
      end
      12'b000101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_365;
      end
      12'b000101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_366;
      end
      12'b000101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_367;
      end
      12'b000101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_368;
      end
      12'b000101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_369;
      end
      12'b000101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_370;
      end
      12'b000101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_371;
      end
      12'b000101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_372;
      end
      12'b000101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_373;
      end
      12'b000101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_374;
      end
      12'b000101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_375;
      end
      12'b000101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_376;
      end
      12'b000101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_377;
      end
      12'b000101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_378;
      end
      12'b000101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_379;
      end
      12'b000101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_380;
      end
      12'b000101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_381;
      end
      12'b000101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_382;
      end
      12'b000101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_383;
      end
      12'b000110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_384;
      end
      12'b000110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_385;
      end
      12'b000110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_386;
      end
      12'b000110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_387;
      end
      12'b000110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_388;
      end
      12'b000110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_389;
      end
      12'b000110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_390;
      end
      12'b000110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_391;
      end
      12'b000110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_392;
      end
      12'b000110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_393;
      end
      12'b000110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_394;
      end
      12'b000110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_395;
      end
      12'b000110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_396;
      end
      12'b000110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_397;
      end
      12'b000110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_398;
      end
      12'b000110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_399;
      end
      12'b000110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_400;
      end
      12'b000110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_401;
      end
      12'b000110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_402;
      end
      12'b000110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_403;
      end
      12'b000110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_404;
      end
      12'b000110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_405;
      end
      12'b000110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_406;
      end
      12'b000110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_407;
      end
      12'b000110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_408;
      end
      12'b000110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_409;
      end
      12'b000110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_410;
      end
      12'b000110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_411;
      end
      12'b000110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_412;
      end
      12'b000110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_413;
      end
      12'b000110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_414;
      end
      12'b000110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_415;
      end
      12'b000110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_416;
      end
      12'b000110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_417;
      end
      12'b000110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_418;
      end
      12'b000110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_419;
      end
      12'b000110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_420;
      end
      12'b000110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_421;
      end
      12'b000110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_422;
      end
      12'b000110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_423;
      end
      12'b000110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_424;
      end
      12'b000110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_425;
      end
      12'b000110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_426;
      end
      12'b000110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_427;
      end
      12'b000110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_428;
      end
      12'b000110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_429;
      end
      12'b000110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_430;
      end
      12'b000110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_431;
      end
      12'b000110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_432;
      end
      12'b000110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_433;
      end
      12'b000110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_434;
      end
      12'b000110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_435;
      end
      12'b000110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_436;
      end
      12'b000110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_437;
      end
      12'b000110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_438;
      end
      12'b000110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_439;
      end
      12'b000110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_440;
      end
      12'b000110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_441;
      end
      12'b000110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_442;
      end
      12'b000110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_443;
      end
      12'b000110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_444;
      end
      12'b000110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_445;
      end
      12'b000110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_446;
      end
      12'b000110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_447;
      end
      12'b000111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_448;
      end
      12'b000111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_449;
      end
      12'b000111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_450;
      end
      12'b000111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_451;
      end
      12'b000111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_452;
      end
      12'b000111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_453;
      end
      12'b000111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_454;
      end
      12'b000111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_455;
      end
      12'b000111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_456;
      end
      12'b000111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_457;
      end
      12'b000111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_458;
      end
      12'b000111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_459;
      end
      12'b000111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_460;
      end
      12'b000111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_461;
      end
      12'b000111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_462;
      end
      12'b000111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_463;
      end
      12'b000111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_464;
      end
      12'b000111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_465;
      end
      12'b000111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_466;
      end
      12'b000111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_467;
      end
      12'b000111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_468;
      end
      12'b000111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_469;
      end
      12'b000111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_470;
      end
      12'b000111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_471;
      end
      12'b000111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_472;
      end
      12'b000111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_473;
      end
      12'b000111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_474;
      end
      12'b000111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_475;
      end
      12'b000111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_476;
      end
      12'b000111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_477;
      end
      12'b000111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_478;
      end
      12'b000111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_479;
      end
      12'b000111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_480;
      end
      12'b000111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_481;
      end
      12'b000111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_482;
      end
      12'b000111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_483;
      end
      12'b000111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_484;
      end
      12'b000111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_485;
      end
      12'b000111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_486;
      end
      12'b000111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_487;
      end
      12'b000111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_488;
      end
      12'b000111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_489;
      end
      12'b000111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_490;
      end
      12'b000111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_491;
      end
      12'b000111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_492;
      end
      12'b000111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_493;
      end
      12'b000111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_494;
      end
      12'b000111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_495;
      end
      12'b000111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_496;
      end
      12'b000111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_497;
      end
      12'b000111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_498;
      end
      12'b000111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_499;
      end
      12'b000111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_500;
      end
      12'b000111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_501;
      end
      12'b000111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_502;
      end
      12'b000111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_503;
      end
      12'b000111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_504;
      end
      12'b000111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_505;
      end
      12'b000111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_506;
      end
      12'b000111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_507;
      end
      12'b000111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_508;
      end
      12'b000111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_509;
      end
      12'b000111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_510;
      end
      12'b000111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_511;
      end
      12'b001000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_512;
      end
      12'b001000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_513;
      end
      12'b001000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_514;
      end
      12'b001000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_515;
      end
      12'b001000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_516;
      end
      12'b001000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_517;
      end
      12'b001000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_518;
      end
      12'b001000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_519;
      end
      12'b001000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_520;
      end
      12'b001000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_521;
      end
      12'b001000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_522;
      end
      12'b001000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_523;
      end
      12'b001000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_524;
      end
      12'b001000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_525;
      end
      12'b001000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_526;
      end
      12'b001000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_527;
      end
      12'b001000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_528;
      end
      12'b001000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_529;
      end
      12'b001000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_530;
      end
      12'b001000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_531;
      end
      12'b001000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_532;
      end
      12'b001000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_533;
      end
      12'b001000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_534;
      end
      12'b001000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_535;
      end
      12'b001000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_536;
      end
      12'b001000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_537;
      end
      12'b001000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_538;
      end
      12'b001000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_539;
      end
      12'b001000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_540;
      end
      12'b001000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_541;
      end
      12'b001000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_542;
      end
      12'b001000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_543;
      end
      12'b001000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_544;
      end
      12'b001000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_545;
      end
      12'b001000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_546;
      end
      12'b001000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_547;
      end
      12'b001000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_548;
      end
      12'b001000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_549;
      end
      12'b001000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_550;
      end
      12'b001000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_551;
      end
      12'b001000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_552;
      end
      12'b001000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_553;
      end
      12'b001000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_554;
      end
      12'b001000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_555;
      end
      12'b001000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_556;
      end
      12'b001000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_557;
      end
      12'b001000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_558;
      end
      12'b001000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_559;
      end
      12'b001000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_560;
      end
      12'b001000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_561;
      end
      12'b001000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_562;
      end
      12'b001000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_563;
      end
      12'b001000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_564;
      end
      12'b001000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_565;
      end
      12'b001000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_566;
      end
      12'b001000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_567;
      end
      12'b001000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_568;
      end
      12'b001000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_569;
      end
      12'b001000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_570;
      end
      12'b001000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_571;
      end
      12'b001000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_572;
      end
      12'b001000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_573;
      end
      12'b001000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_574;
      end
      12'b001000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_575;
      end
      12'b001001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_576;
      end
      12'b001001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_577;
      end
      12'b001001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_578;
      end
      12'b001001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_579;
      end
      12'b001001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_580;
      end
      12'b001001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_581;
      end
      12'b001001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_582;
      end
      12'b001001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_583;
      end
      12'b001001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_584;
      end
      12'b001001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_585;
      end
      12'b001001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_586;
      end
      12'b001001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_587;
      end
      12'b001001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_588;
      end
      12'b001001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_589;
      end
      12'b001001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_590;
      end
      12'b001001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_591;
      end
      12'b001001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_592;
      end
      12'b001001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_593;
      end
      12'b001001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_594;
      end
      12'b001001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_595;
      end
      12'b001001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_596;
      end
      12'b001001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_597;
      end
      12'b001001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_598;
      end
      12'b001001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_599;
      end
      12'b001001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_600;
      end
      12'b001001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_601;
      end
      12'b001001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_602;
      end
      12'b001001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_603;
      end
      12'b001001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_604;
      end
      12'b001001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_605;
      end
      12'b001001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_606;
      end
      12'b001001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_607;
      end
      12'b001001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_608;
      end
      12'b001001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_609;
      end
      12'b001001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_610;
      end
      12'b001001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_611;
      end
      12'b001001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_612;
      end
      12'b001001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_613;
      end
      12'b001001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_614;
      end
      12'b001001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_615;
      end
      12'b001001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_616;
      end
      12'b001001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_617;
      end
      12'b001001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_618;
      end
      12'b001001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_619;
      end
      12'b001001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_620;
      end
      12'b001001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_621;
      end
      12'b001001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_622;
      end
      12'b001001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_623;
      end
      12'b001001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_624;
      end
      12'b001001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_625;
      end
      12'b001001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_626;
      end
      12'b001001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_627;
      end
      12'b001001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_628;
      end
      12'b001001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_629;
      end
      12'b001001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_630;
      end
      12'b001001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_631;
      end
      12'b001001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_632;
      end
      12'b001001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_633;
      end
      12'b001001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_634;
      end
      12'b001001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_635;
      end
      12'b001001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_636;
      end
      12'b001001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_637;
      end
      12'b001001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_638;
      end
      12'b001001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_639;
      end
      12'b001010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_640;
      end
      12'b001010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_641;
      end
      12'b001010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_642;
      end
      12'b001010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_643;
      end
      12'b001010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_644;
      end
      12'b001010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_645;
      end
      12'b001010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_646;
      end
      12'b001010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_647;
      end
      12'b001010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_648;
      end
      12'b001010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_649;
      end
      12'b001010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_650;
      end
      12'b001010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_651;
      end
      12'b001010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_652;
      end
      12'b001010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_653;
      end
      12'b001010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_654;
      end
      12'b001010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_655;
      end
      12'b001010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_656;
      end
      12'b001010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_657;
      end
      12'b001010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_658;
      end
      12'b001010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_659;
      end
      12'b001010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_660;
      end
      12'b001010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_661;
      end
      12'b001010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_662;
      end
      12'b001010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_663;
      end
      12'b001010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_664;
      end
      12'b001010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_665;
      end
      12'b001010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_666;
      end
      12'b001010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_667;
      end
      12'b001010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_668;
      end
      12'b001010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_669;
      end
      12'b001010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_670;
      end
      12'b001010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_671;
      end
      12'b001010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_672;
      end
      12'b001010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_673;
      end
      12'b001010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_674;
      end
      12'b001010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_675;
      end
      12'b001010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_676;
      end
      12'b001010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_677;
      end
      12'b001010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_678;
      end
      12'b001010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_679;
      end
      12'b001010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_680;
      end
      12'b001010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_681;
      end
      12'b001010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_682;
      end
      12'b001010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_683;
      end
      12'b001010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_684;
      end
      12'b001010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_685;
      end
      12'b001010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_686;
      end
      12'b001010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_687;
      end
      12'b001010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_688;
      end
      12'b001010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_689;
      end
      12'b001010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_690;
      end
      12'b001010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_691;
      end
      12'b001010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_692;
      end
      12'b001010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_693;
      end
      12'b001010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_694;
      end
      12'b001010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_695;
      end
      12'b001010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_696;
      end
      12'b001010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_697;
      end
      12'b001010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_698;
      end
      12'b001010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_699;
      end
      12'b001010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_700;
      end
      12'b001010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_701;
      end
      12'b001010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_702;
      end
      12'b001010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_703;
      end
      12'b001011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_704;
      end
      12'b001011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_705;
      end
      12'b001011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_706;
      end
      12'b001011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_707;
      end
      12'b001011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_708;
      end
      12'b001011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_709;
      end
      12'b001011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_710;
      end
      12'b001011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_711;
      end
      12'b001011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_712;
      end
      12'b001011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_713;
      end
      12'b001011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_714;
      end
      12'b001011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_715;
      end
      12'b001011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_716;
      end
      12'b001011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_717;
      end
      12'b001011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_718;
      end
      12'b001011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_719;
      end
      12'b001011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_720;
      end
      12'b001011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_721;
      end
      12'b001011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_722;
      end
      12'b001011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_723;
      end
      12'b001011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_724;
      end
      12'b001011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_725;
      end
      12'b001011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_726;
      end
      12'b001011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_727;
      end
      12'b001011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_728;
      end
      12'b001011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_729;
      end
      12'b001011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_730;
      end
      12'b001011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_731;
      end
      12'b001011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_732;
      end
      12'b001011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_733;
      end
      12'b001011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_734;
      end
      12'b001011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_735;
      end
      12'b001011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_736;
      end
      12'b001011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_737;
      end
      12'b001011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_738;
      end
      12'b001011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_739;
      end
      12'b001011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_740;
      end
      12'b001011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_741;
      end
      12'b001011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_742;
      end
      12'b001011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_743;
      end
      12'b001011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_744;
      end
      12'b001011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_745;
      end
      12'b001011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_746;
      end
      12'b001011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_747;
      end
      12'b001011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_748;
      end
      12'b001011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_749;
      end
      12'b001011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_750;
      end
      12'b001011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_751;
      end
      12'b001011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_752;
      end
      12'b001011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_753;
      end
      12'b001011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_754;
      end
      12'b001011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_755;
      end
      12'b001011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_756;
      end
      12'b001011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_757;
      end
      12'b001011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_758;
      end
      12'b001011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_759;
      end
      12'b001011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_760;
      end
      12'b001011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_761;
      end
      12'b001011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_762;
      end
      12'b001011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_763;
      end
      12'b001011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_764;
      end
      12'b001011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_765;
      end
      12'b001011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_766;
      end
      12'b001011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_767;
      end
      12'b001100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_768;
      end
      12'b001100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_769;
      end
      12'b001100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_770;
      end
      12'b001100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_771;
      end
      12'b001100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_772;
      end
      12'b001100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_773;
      end
      12'b001100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_774;
      end
      12'b001100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_775;
      end
      12'b001100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_776;
      end
      12'b001100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_777;
      end
      12'b001100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_778;
      end
      12'b001100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_779;
      end
      12'b001100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_780;
      end
      12'b001100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_781;
      end
      12'b001100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_782;
      end
      12'b001100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_783;
      end
      12'b001100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_784;
      end
      12'b001100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_785;
      end
      12'b001100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_786;
      end
      12'b001100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_787;
      end
      12'b001100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_788;
      end
      12'b001100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_789;
      end
      12'b001100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_790;
      end
      12'b001100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_791;
      end
      12'b001100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_792;
      end
      12'b001100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_793;
      end
      12'b001100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_794;
      end
      12'b001100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_795;
      end
      12'b001100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_796;
      end
      12'b001100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_797;
      end
      12'b001100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_798;
      end
      12'b001100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_799;
      end
      12'b001100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_800;
      end
      12'b001100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_801;
      end
      12'b001100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_802;
      end
      12'b001100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_803;
      end
      12'b001100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_804;
      end
      12'b001100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_805;
      end
      12'b001100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_806;
      end
      12'b001100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_807;
      end
      12'b001100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_808;
      end
      12'b001100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_809;
      end
      12'b001100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_810;
      end
      12'b001100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_811;
      end
      12'b001100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_812;
      end
      12'b001100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_813;
      end
      12'b001100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_814;
      end
      12'b001100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_815;
      end
      12'b001100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_816;
      end
      12'b001100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_817;
      end
      12'b001100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_818;
      end
      12'b001100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_819;
      end
      12'b001100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_820;
      end
      12'b001100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_821;
      end
      12'b001100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_822;
      end
      12'b001100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_823;
      end
      12'b001100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_824;
      end
      12'b001100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_825;
      end
      12'b001100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_826;
      end
      12'b001100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_827;
      end
      12'b001100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_828;
      end
      12'b001100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_829;
      end
      12'b001100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_830;
      end
      12'b001100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_831;
      end
      12'b001101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_832;
      end
      12'b001101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_833;
      end
      12'b001101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_834;
      end
      12'b001101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_835;
      end
      12'b001101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_836;
      end
      12'b001101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_837;
      end
      12'b001101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_838;
      end
      12'b001101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_839;
      end
      12'b001101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_840;
      end
      12'b001101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_841;
      end
      12'b001101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_842;
      end
      12'b001101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_843;
      end
      12'b001101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_844;
      end
      12'b001101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_845;
      end
      12'b001101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_846;
      end
      12'b001101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_847;
      end
      12'b001101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_848;
      end
      12'b001101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_849;
      end
      12'b001101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_850;
      end
      12'b001101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_851;
      end
      12'b001101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_852;
      end
      12'b001101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_853;
      end
      12'b001101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_854;
      end
      12'b001101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_855;
      end
      12'b001101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_856;
      end
      12'b001101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_857;
      end
      12'b001101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_858;
      end
      12'b001101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_859;
      end
      12'b001101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_860;
      end
      12'b001101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_861;
      end
      12'b001101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_862;
      end
      12'b001101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_863;
      end
      12'b001101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_864;
      end
      12'b001101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_865;
      end
      12'b001101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_866;
      end
      12'b001101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_867;
      end
      12'b001101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_868;
      end
      12'b001101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_869;
      end
      12'b001101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_870;
      end
      12'b001101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_871;
      end
      12'b001101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_872;
      end
      12'b001101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_873;
      end
      12'b001101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_874;
      end
      12'b001101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_875;
      end
      12'b001101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_876;
      end
      12'b001101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_877;
      end
      12'b001101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_878;
      end
      12'b001101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_879;
      end
      12'b001101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_880;
      end
      12'b001101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_881;
      end
      12'b001101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_882;
      end
      12'b001101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_883;
      end
      12'b001101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_884;
      end
      12'b001101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_885;
      end
      12'b001101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_886;
      end
      12'b001101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_887;
      end
      12'b001101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_888;
      end
      12'b001101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_889;
      end
      12'b001101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_890;
      end
      12'b001101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_891;
      end
      12'b001101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_892;
      end
      12'b001101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_893;
      end
      12'b001101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_894;
      end
      12'b001101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_895;
      end
      12'b001110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_896;
      end
      12'b001110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_897;
      end
      12'b001110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_898;
      end
      12'b001110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_899;
      end
      12'b001110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_900;
      end
      12'b001110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_901;
      end
      12'b001110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_902;
      end
      12'b001110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_903;
      end
      12'b001110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_904;
      end
      12'b001110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_905;
      end
      12'b001110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_906;
      end
      12'b001110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_907;
      end
      12'b001110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_908;
      end
      12'b001110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_909;
      end
      12'b001110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_910;
      end
      12'b001110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_911;
      end
      12'b001110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_912;
      end
      12'b001110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_913;
      end
      12'b001110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_914;
      end
      12'b001110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_915;
      end
      12'b001110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_916;
      end
      12'b001110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_917;
      end
      12'b001110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_918;
      end
      12'b001110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_919;
      end
      12'b001110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_920;
      end
      12'b001110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_921;
      end
      12'b001110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_922;
      end
      12'b001110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_923;
      end
      12'b001110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_924;
      end
      12'b001110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_925;
      end
      12'b001110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_926;
      end
      12'b001110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_927;
      end
      12'b001110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_928;
      end
      12'b001110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_929;
      end
      12'b001110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_930;
      end
      12'b001110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_931;
      end
      12'b001110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_932;
      end
      12'b001110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_933;
      end
      12'b001110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_934;
      end
      12'b001110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_935;
      end
      12'b001110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_936;
      end
      12'b001110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_937;
      end
      12'b001110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_938;
      end
      12'b001110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_939;
      end
      12'b001110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_940;
      end
      12'b001110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_941;
      end
      12'b001110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_942;
      end
      12'b001110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_943;
      end
      12'b001110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_944;
      end
      12'b001110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_945;
      end
      12'b001110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_946;
      end
      12'b001110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_947;
      end
      12'b001110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_948;
      end
      12'b001110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_949;
      end
      12'b001110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_950;
      end
      12'b001110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_951;
      end
      12'b001110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_952;
      end
      12'b001110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_953;
      end
      12'b001110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_954;
      end
      12'b001110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_955;
      end
      12'b001110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_956;
      end
      12'b001110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_957;
      end
      12'b001110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_958;
      end
      12'b001110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_959;
      end
      12'b001111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_960;
      end
      12'b001111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_961;
      end
      12'b001111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_962;
      end
      12'b001111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_963;
      end
      12'b001111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_964;
      end
      12'b001111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_965;
      end
      12'b001111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_966;
      end
      12'b001111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_967;
      end
      12'b001111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_968;
      end
      12'b001111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_969;
      end
      12'b001111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_970;
      end
      12'b001111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_971;
      end
      12'b001111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_972;
      end
      12'b001111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_973;
      end
      12'b001111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_974;
      end
      12'b001111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_975;
      end
      12'b001111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_976;
      end
      12'b001111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_977;
      end
      12'b001111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_978;
      end
      12'b001111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_979;
      end
      12'b001111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_980;
      end
      12'b001111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_981;
      end
      12'b001111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_982;
      end
      12'b001111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_983;
      end
      12'b001111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_984;
      end
      12'b001111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_985;
      end
      12'b001111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_986;
      end
      12'b001111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_987;
      end
      12'b001111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_988;
      end
      12'b001111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_989;
      end
      12'b001111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_990;
      end
      12'b001111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_991;
      end
      12'b001111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_992;
      end
      12'b001111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_993;
      end
      12'b001111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_994;
      end
      12'b001111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_995;
      end
      12'b001111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_996;
      end
      12'b001111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_997;
      end
      12'b001111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_998;
      end
      12'b001111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_999;
      end
      12'b001111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1000;
      end
      12'b001111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1001;
      end
      12'b001111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1002;
      end
      12'b001111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1003;
      end
      12'b001111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1004;
      end
      12'b001111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1005;
      end
      12'b001111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1006;
      end
      12'b001111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1007;
      end
      12'b001111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1008;
      end
      12'b001111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1009;
      end
      12'b001111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1010;
      end
      12'b001111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1011;
      end
      12'b001111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1012;
      end
      12'b001111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1013;
      end
      12'b001111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1014;
      end
      12'b001111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1015;
      end
      12'b001111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1016;
      end
      12'b001111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1017;
      end
      12'b001111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1018;
      end
      12'b001111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1019;
      end
      12'b001111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1020;
      end
      12'b001111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1021;
      end
      12'b001111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1022;
      end
      12'b001111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1023;
      end
      12'b010000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1024;
      end
      12'b010000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1025;
      end
      12'b010000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1026;
      end
      12'b010000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1027;
      end
      12'b010000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1028;
      end
      12'b010000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1029;
      end
      12'b010000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1030;
      end
      12'b010000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1031;
      end
      12'b010000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1032;
      end
      12'b010000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1033;
      end
      12'b010000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1034;
      end
      12'b010000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1035;
      end
      12'b010000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1036;
      end
      12'b010000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1037;
      end
      12'b010000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1038;
      end
      12'b010000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1039;
      end
      12'b010000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1040;
      end
      12'b010000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1041;
      end
      12'b010000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1042;
      end
      12'b010000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1043;
      end
      12'b010000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1044;
      end
      12'b010000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1045;
      end
      12'b010000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1046;
      end
      12'b010000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1047;
      end
      12'b010000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1048;
      end
      12'b010000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1049;
      end
      12'b010000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1050;
      end
      12'b010000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1051;
      end
      12'b010000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1052;
      end
      12'b010000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1053;
      end
      12'b010000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1054;
      end
      12'b010000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1055;
      end
      12'b010000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1056;
      end
      12'b010000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1057;
      end
      12'b010000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1058;
      end
      12'b010000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1059;
      end
      12'b010000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1060;
      end
      12'b010000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1061;
      end
      12'b010000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1062;
      end
      12'b010000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1063;
      end
      12'b010000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1064;
      end
      12'b010000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1065;
      end
      12'b010000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1066;
      end
      12'b010000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1067;
      end
      12'b010000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1068;
      end
      12'b010000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1069;
      end
      12'b010000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1070;
      end
      12'b010000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1071;
      end
      12'b010000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1072;
      end
      12'b010000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1073;
      end
      12'b010000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1074;
      end
      12'b010000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1075;
      end
      12'b010000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1076;
      end
      12'b010000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1077;
      end
      12'b010000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1078;
      end
      12'b010000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1079;
      end
      12'b010000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1080;
      end
      12'b010000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1081;
      end
      12'b010000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1082;
      end
      12'b010000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1083;
      end
      12'b010000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1084;
      end
      12'b010000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1085;
      end
      12'b010000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1086;
      end
      12'b010000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1087;
      end
      12'b010001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1088;
      end
      12'b010001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1089;
      end
      12'b010001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1090;
      end
      12'b010001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1091;
      end
      12'b010001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1092;
      end
      12'b010001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1093;
      end
      12'b010001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1094;
      end
      12'b010001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1095;
      end
      12'b010001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1096;
      end
      12'b010001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1097;
      end
      12'b010001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1098;
      end
      12'b010001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1099;
      end
      12'b010001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1100;
      end
      12'b010001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1101;
      end
      12'b010001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1102;
      end
      12'b010001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1103;
      end
      12'b010001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1104;
      end
      12'b010001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1105;
      end
      12'b010001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1106;
      end
      12'b010001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1107;
      end
      12'b010001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1108;
      end
      12'b010001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1109;
      end
      12'b010001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1110;
      end
      12'b010001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1111;
      end
      12'b010001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1112;
      end
      12'b010001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1113;
      end
      12'b010001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1114;
      end
      12'b010001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1115;
      end
      12'b010001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1116;
      end
      12'b010001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1117;
      end
      12'b010001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1118;
      end
      12'b010001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1119;
      end
      12'b010001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1120;
      end
      12'b010001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1121;
      end
      12'b010001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1122;
      end
      12'b010001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1123;
      end
      12'b010001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1124;
      end
      12'b010001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1125;
      end
      12'b010001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1126;
      end
      12'b010001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1127;
      end
      12'b010001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1128;
      end
      12'b010001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1129;
      end
      12'b010001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1130;
      end
      12'b010001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1131;
      end
      12'b010001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1132;
      end
      12'b010001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1133;
      end
      12'b010001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1134;
      end
      12'b010001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1135;
      end
      12'b010001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1136;
      end
      12'b010001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1137;
      end
      12'b010001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1138;
      end
      12'b010001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1139;
      end
      12'b010001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1140;
      end
      12'b010001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1141;
      end
      12'b010001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1142;
      end
      12'b010001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1143;
      end
      12'b010001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1144;
      end
      12'b010001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1145;
      end
      12'b010001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1146;
      end
      12'b010001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1147;
      end
      12'b010001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1148;
      end
      12'b010001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1149;
      end
      12'b010001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1150;
      end
      12'b010001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1151;
      end
      12'b010010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1152;
      end
      12'b010010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1153;
      end
      12'b010010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1154;
      end
      12'b010010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1155;
      end
      12'b010010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1156;
      end
      12'b010010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1157;
      end
      12'b010010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1158;
      end
      12'b010010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1159;
      end
      12'b010010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1160;
      end
      12'b010010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1161;
      end
      12'b010010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1162;
      end
      12'b010010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1163;
      end
      12'b010010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1164;
      end
      12'b010010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1165;
      end
      12'b010010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1166;
      end
      12'b010010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1167;
      end
      12'b010010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1168;
      end
      12'b010010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1169;
      end
      12'b010010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1170;
      end
      12'b010010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1171;
      end
      12'b010010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1172;
      end
      12'b010010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1173;
      end
      12'b010010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1174;
      end
      12'b010010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1175;
      end
      12'b010010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1176;
      end
      12'b010010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1177;
      end
      12'b010010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1178;
      end
      12'b010010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1179;
      end
      12'b010010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1180;
      end
      12'b010010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1181;
      end
      12'b010010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1182;
      end
      12'b010010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1183;
      end
      12'b010010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1184;
      end
      12'b010010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1185;
      end
      12'b010010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1186;
      end
      12'b010010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1187;
      end
      12'b010010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1188;
      end
      12'b010010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1189;
      end
      12'b010010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1190;
      end
      12'b010010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1191;
      end
      12'b010010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1192;
      end
      12'b010010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1193;
      end
      12'b010010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1194;
      end
      12'b010010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1195;
      end
      12'b010010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1196;
      end
      12'b010010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1197;
      end
      12'b010010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1198;
      end
      12'b010010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1199;
      end
      12'b010010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1200;
      end
      12'b010010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1201;
      end
      12'b010010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1202;
      end
      12'b010010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1203;
      end
      12'b010010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1204;
      end
      12'b010010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1205;
      end
      12'b010010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1206;
      end
      12'b010010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1207;
      end
      12'b010010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1208;
      end
      12'b010010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1209;
      end
      12'b010010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1210;
      end
      12'b010010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1211;
      end
      12'b010010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1212;
      end
      12'b010010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1213;
      end
      12'b010010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1214;
      end
      12'b010010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1215;
      end
      12'b010011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1216;
      end
      12'b010011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1217;
      end
      12'b010011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1218;
      end
      12'b010011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1219;
      end
      12'b010011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1220;
      end
      12'b010011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1221;
      end
      12'b010011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1222;
      end
      12'b010011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1223;
      end
      12'b010011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1224;
      end
      12'b010011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1225;
      end
      12'b010011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1226;
      end
      12'b010011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1227;
      end
      12'b010011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1228;
      end
      12'b010011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1229;
      end
      12'b010011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1230;
      end
      12'b010011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1231;
      end
      12'b010011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1232;
      end
      12'b010011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1233;
      end
      12'b010011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1234;
      end
      12'b010011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1235;
      end
      12'b010011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1236;
      end
      12'b010011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1237;
      end
      12'b010011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1238;
      end
      12'b010011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1239;
      end
      12'b010011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1240;
      end
      12'b010011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1241;
      end
      12'b010011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1242;
      end
      12'b010011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1243;
      end
      12'b010011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1244;
      end
      12'b010011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1245;
      end
      12'b010011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1246;
      end
      12'b010011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1247;
      end
      12'b010011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1248;
      end
      12'b010011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1249;
      end
      12'b010011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1250;
      end
      12'b010011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1251;
      end
      12'b010011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1252;
      end
      12'b010011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1253;
      end
      12'b010011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1254;
      end
      12'b010011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1255;
      end
      12'b010011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1256;
      end
      12'b010011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1257;
      end
      12'b010011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1258;
      end
      12'b010011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1259;
      end
      12'b010011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1260;
      end
      12'b010011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1261;
      end
      12'b010011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1262;
      end
      12'b010011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1263;
      end
      12'b010011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1264;
      end
      12'b010011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1265;
      end
      12'b010011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1266;
      end
      12'b010011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1267;
      end
      12'b010011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1268;
      end
      12'b010011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1269;
      end
      12'b010011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1270;
      end
      12'b010011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1271;
      end
      12'b010011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1272;
      end
      12'b010011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1273;
      end
      12'b010011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1274;
      end
      12'b010011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1275;
      end
      12'b010011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1276;
      end
      12'b010011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1277;
      end
      12'b010011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1278;
      end
      12'b010011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1279;
      end
      12'b010100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1280;
      end
      12'b010100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1281;
      end
      12'b010100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1282;
      end
      12'b010100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1283;
      end
      12'b010100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1284;
      end
      12'b010100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1285;
      end
      12'b010100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1286;
      end
      12'b010100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1287;
      end
      12'b010100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1288;
      end
      12'b010100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1289;
      end
      12'b010100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1290;
      end
      12'b010100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1291;
      end
      12'b010100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1292;
      end
      12'b010100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1293;
      end
      12'b010100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1294;
      end
      12'b010100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1295;
      end
      12'b010100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1296;
      end
      12'b010100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1297;
      end
      12'b010100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1298;
      end
      12'b010100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1299;
      end
      12'b010100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1300;
      end
      12'b010100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1301;
      end
      12'b010100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1302;
      end
      12'b010100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1303;
      end
      12'b010100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1304;
      end
      12'b010100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1305;
      end
      12'b010100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1306;
      end
      12'b010100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1307;
      end
      12'b010100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1308;
      end
      12'b010100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1309;
      end
      12'b010100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1310;
      end
      12'b010100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1311;
      end
      12'b010100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1312;
      end
      12'b010100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1313;
      end
      12'b010100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1314;
      end
      12'b010100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1315;
      end
      12'b010100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1316;
      end
      12'b010100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1317;
      end
      12'b010100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1318;
      end
      12'b010100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1319;
      end
      12'b010100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1320;
      end
      12'b010100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1321;
      end
      12'b010100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1322;
      end
      12'b010100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1323;
      end
      12'b010100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1324;
      end
      12'b010100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1325;
      end
      12'b010100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1326;
      end
      12'b010100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1327;
      end
      12'b010100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1328;
      end
      12'b010100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1329;
      end
      12'b010100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1330;
      end
      12'b010100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1331;
      end
      12'b010100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1332;
      end
      12'b010100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1333;
      end
      12'b010100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1334;
      end
      12'b010100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1335;
      end
      12'b010100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1336;
      end
      12'b010100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1337;
      end
      12'b010100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1338;
      end
      12'b010100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1339;
      end
      12'b010100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1340;
      end
      12'b010100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1341;
      end
      12'b010100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1342;
      end
      12'b010100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1343;
      end
      12'b010101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1344;
      end
      12'b010101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1345;
      end
      12'b010101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1346;
      end
      12'b010101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1347;
      end
      12'b010101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1348;
      end
      12'b010101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1349;
      end
      12'b010101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1350;
      end
      12'b010101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1351;
      end
      12'b010101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1352;
      end
      12'b010101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1353;
      end
      12'b010101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1354;
      end
      12'b010101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1355;
      end
      12'b010101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1356;
      end
      12'b010101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1357;
      end
      12'b010101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1358;
      end
      12'b010101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1359;
      end
      12'b010101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1360;
      end
      12'b010101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1361;
      end
      12'b010101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1362;
      end
      12'b010101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1363;
      end
      12'b010101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1364;
      end
      12'b010101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1365;
      end
      12'b010101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1366;
      end
      12'b010101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1367;
      end
      12'b010101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1368;
      end
      12'b010101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1369;
      end
      12'b010101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1370;
      end
      12'b010101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1371;
      end
      12'b010101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1372;
      end
      12'b010101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1373;
      end
      12'b010101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1374;
      end
      12'b010101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1375;
      end
      12'b010101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1376;
      end
      12'b010101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1377;
      end
      12'b010101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1378;
      end
      12'b010101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1379;
      end
      12'b010101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1380;
      end
      12'b010101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1381;
      end
      12'b010101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1382;
      end
      12'b010101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1383;
      end
      12'b010101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1384;
      end
      12'b010101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1385;
      end
      12'b010101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1386;
      end
      12'b010101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1387;
      end
      12'b010101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1388;
      end
      12'b010101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1389;
      end
      12'b010101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1390;
      end
      12'b010101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1391;
      end
      12'b010101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1392;
      end
      12'b010101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1393;
      end
      12'b010101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1394;
      end
      12'b010101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1395;
      end
      12'b010101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1396;
      end
      12'b010101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1397;
      end
      12'b010101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1398;
      end
      12'b010101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1399;
      end
      12'b010101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1400;
      end
      12'b010101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1401;
      end
      12'b010101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1402;
      end
      12'b010101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1403;
      end
      12'b010101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1404;
      end
      12'b010101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1405;
      end
      12'b010101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1406;
      end
      12'b010101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1407;
      end
      12'b010110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1408;
      end
      12'b010110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1409;
      end
      12'b010110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1410;
      end
      12'b010110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1411;
      end
      12'b010110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1412;
      end
      12'b010110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1413;
      end
      12'b010110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1414;
      end
      12'b010110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1415;
      end
      12'b010110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1416;
      end
      12'b010110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1417;
      end
      12'b010110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1418;
      end
      12'b010110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1419;
      end
      12'b010110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1420;
      end
      12'b010110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1421;
      end
      12'b010110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1422;
      end
      12'b010110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1423;
      end
      12'b010110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1424;
      end
      12'b010110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1425;
      end
      12'b010110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1426;
      end
      12'b010110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1427;
      end
      12'b010110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1428;
      end
      12'b010110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1429;
      end
      12'b010110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1430;
      end
      12'b010110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1431;
      end
      12'b010110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1432;
      end
      12'b010110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1433;
      end
      12'b010110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1434;
      end
      12'b010110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1435;
      end
      12'b010110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1436;
      end
      12'b010110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1437;
      end
      12'b010110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1438;
      end
      12'b010110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1439;
      end
      12'b010110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1440;
      end
      12'b010110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1441;
      end
      12'b010110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1442;
      end
      12'b010110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1443;
      end
      12'b010110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1444;
      end
      12'b010110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1445;
      end
      12'b010110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1446;
      end
      12'b010110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1447;
      end
      12'b010110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1448;
      end
      12'b010110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1449;
      end
      12'b010110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1450;
      end
      12'b010110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1451;
      end
      12'b010110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1452;
      end
      12'b010110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1453;
      end
      12'b010110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1454;
      end
      12'b010110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1455;
      end
      12'b010110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1456;
      end
      12'b010110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1457;
      end
      12'b010110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1458;
      end
      12'b010110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1459;
      end
      12'b010110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1460;
      end
      12'b010110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1461;
      end
      12'b010110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1462;
      end
      12'b010110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1463;
      end
      12'b010110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1464;
      end
      12'b010110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1465;
      end
      12'b010110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1466;
      end
      12'b010110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1467;
      end
      12'b010110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1468;
      end
      12'b010110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1469;
      end
      12'b010110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1470;
      end
      12'b010110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1471;
      end
      12'b010111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1472;
      end
      12'b010111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1473;
      end
      12'b010111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1474;
      end
      12'b010111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1475;
      end
      12'b010111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1476;
      end
      12'b010111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1477;
      end
      12'b010111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1478;
      end
      12'b010111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1479;
      end
      12'b010111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1480;
      end
      12'b010111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1481;
      end
      12'b010111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1482;
      end
      12'b010111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1483;
      end
      12'b010111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1484;
      end
      12'b010111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1485;
      end
      12'b010111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1486;
      end
      12'b010111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1487;
      end
      12'b010111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1488;
      end
      12'b010111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1489;
      end
      12'b010111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1490;
      end
      12'b010111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1491;
      end
      12'b010111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1492;
      end
      12'b010111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1493;
      end
      12'b010111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1494;
      end
      12'b010111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1495;
      end
      12'b010111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1496;
      end
      12'b010111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1497;
      end
      12'b010111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1498;
      end
      12'b010111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1499;
      end
      12'b010111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1500;
      end
      12'b010111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1501;
      end
      12'b010111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1502;
      end
      12'b010111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1503;
      end
      12'b010111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1504;
      end
      12'b010111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1505;
      end
      12'b010111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1506;
      end
      12'b010111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1507;
      end
      12'b010111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1508;
      end
      12'b010111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1509;
      end
      12'b010111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1510;
      end
      12'b010111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1511;
      end
      12'b010111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1512;
      end
      12'b010111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1513;
      end
      12'b010111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1514;
      end
      12'b010111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1515;
      end
      12'b010111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1516;
      end
      12'b010111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1517;
      end
      12'b010111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1518;
      end
      12'b010111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1519;
      end
      12'b010111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1520;
      end
      12'b010111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1521;
      end
      12'b010111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1522;
      end
      12'b010111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1523;
      end
      12'b010111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1524;
      end
      12'b010111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1525;
      end
      12'b010111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1526;
      end
      12'b010111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1527;
      end
      12'b010111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1528;
      end
      12'b010111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1529;
      end
      12'b010111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1530;
      end
      12'b010111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1531;
      end
      12'b010111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1532;
      end
      12'b010111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1533;
      end
      12'b010111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1534;
      end
      12'b010111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1535;
      end
      12'b011000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1536;
      end
      12'b011000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1537;
      end
      12'b011000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1538;
      end
      12'b011000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1539;
      end
      12'b011000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1540;
      end
      12'b011000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1541;
      end
      12'b011000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1542;
      end
      12'b011000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1543;
      end
      12'b011000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1544;
      end
      12'b011000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1545;
      end
      12'b011000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1546;
      end
      12'b011000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1547;
      end
      12'b011000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1548;
      end
      12'b011000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1549;
      end
      12'b011000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1550;
      end
      12'b011000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1551;
      end
      12'b011000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1552;
      end
      12'b011000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1553;
      end
      12'b011000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1554;
      end
      12'b011000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1555;
      end
      12'b011000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1556;
      end
      12'b011000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1557;
      end
      12'b011000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1558;
      end
      12'b011000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1559;
      end
      12'b011000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1560;
      end
      12'b011000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1561;
      end
      12'b011000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1562;
      end
      12'b011000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1563;
      end
      12'b011000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1564;
      end
      12'b011000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1565;
      end
      12'b011000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1566;
      end
      12'b011000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1567;
      end
      12'b011000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1568;
      end
      12'b011000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1569;
      end
      12'b011000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1570;
      end
      12'b011000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1571;
      end
      12'b011000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1572;
      end
      12'b011000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1573;
      end
      12'b011000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1574;
      end
      12'b011000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1575;
      end
      12'b011000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1576;
      end
      12'b011000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1577;
      end
      12'b011000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1578;
      end
      12'b011000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1579;
      end
      12'b011000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1580;
      end
      12'b011000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1581;
      end
      12'b011000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1582;
      end
      12'b011000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1583;
      end
      12'b011000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1584;
      end
      12'b011000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1585;
      end
      12'b011000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1586;
      end
      12'b011000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1587;
      end
      12'b011000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1588;
      end
      12'b011000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1589;
      end
      12'b011000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1590;
      end
      12'b011000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1591;
      end
      12'b011000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1592;
      end
      12'b011000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1593;
      end
      12'b011000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1594;
      end
      12'b011000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1595;
      end
      12'b011000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1596;
      end
      12'b011000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1597;
      end
      12'b011000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1598;
      end
      12'b011000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1599;
      end
      12'b011001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1600;
      end
      12'b011001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1601;
      end
      12'b011001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1602;
      end
      12'b011001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1603;
      end
      12'b011001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1604;
      end
      12'b011001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1605;
      end
      12'b011001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1606;
      end
      12'b011001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1607;
      end
      12'b011001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1608;
      end
      12'b011001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1609;
      end
      12'b011001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1610;
      end
      12'b011001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1611;
      end
      12'b011001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1612;
      end
      12'b011001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1613;
      end
      12'b011001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1614;
      end
      12'b011001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1615;
      end
      12'b011001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1616;
      end
      12'b011001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1617;
      end
      12'b011001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1618;
      end
      12'b011001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1619;
      end
      12'b011001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1620;
      end
      12'b011001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1621;
      end
      12'b011001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1622;
      end
      12'b011001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1623;
      end
      12'b011001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1624;
      end
      12'b011001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1625;
      end
      12'b011001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1626;
      end
      12'b011001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1627;
      end
      12'b011001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1628;
      end
      12'b011001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1629;
      end
      12'b011001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1630;
      end
      12'b011001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1631;
      end
      12'b011001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1632;
      end
      12'b011001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1633;
      end
      12'b011001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1634;
      end
      12'b011001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1635;
      end
      12'b011001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1636;
      end
      12'b011001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1637;
      end
      12'b011001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1638;
      end
      12'b011001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1639;
      end
      12'b011001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1640;
      end
      12'b011001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1641;
      end
      12'b011001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1642;
      end
      12'b011001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1643;
      end
      12'b011001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1644;
      end
      12'b011001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1645;
      end
      12'b011001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1646;
      end
      12'b011001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1647;
      end
      12'b011001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1648;
      end
      12'b011001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1649;
      end
      12'b011001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1650;
      end
      12'b011001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1651;
      end
      12'b011001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1652;
      end
      12'b011001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1653;
      end
      12'b011001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1654;
      end
      12'b011001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1655;
      end
      12'b011001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1656;
      end
      12'b011001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1657;
      end
      12'b011001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1658;
      end
      12'b011001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1659;
      end
      12'b011001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1660;
      end
      12'b011001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1661;
      end
      12'b011001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1662;
      end
      12'b011001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1663;
      end
      12'b011010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1664;
      end
      12'b011010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1665;
      end
      12'b011010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1666;
      end
      12'b011010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1667;
      end
      12'b011010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1668;
      end
      12'b011010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1669;
      end
      12'b011010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1670;
      end
      12'b011010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1671;
      end
      12'b011010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1672;
      end
      12'b011010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1673;
      end
      12'b011010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1674;
      end
      12'b011010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1675;
      end
      12'b011010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1676;
      end
      12'b011010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1677;
      end
      12'b011010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1678;
      end
      12'b011010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1679;
      end
      12'b011010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1680;
      end
      12'b011010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1681;
      end
      12'b011010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1682;
      end
      12'b011010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1683;
      end
      12'b011010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1684;
      end
      12'b011010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1685;
      end
      12'b011010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1686;
      end
      12'b011010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1687;
      end
      12'b011010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1688;
      end
      12'b011010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1689;
      end
      12'b011010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1690;
      end
      12'b011010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1691;
      end
      12'b011010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1692;
      end
      12'b011010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1693;
      end
      12'b011010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1694;
      end
      12'b011010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1695;
      end
      12'b011010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1696;
      end
      12'b011010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1697;
      end
      12'b011010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1698;
      end
      12'b011010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1699;
      end
      12'b011010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1700;
      end
      12'b011010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1701;
      end
      12'b011010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1702;
      end
      12'b011010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1703;
      end
      12'b011010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1704;
      end
      12'b011010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1705;
      end
      12'b011010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1706;
      end
      12'b011010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1707;
      end
      12'b011010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1708;
      end
      12'b011010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1709;
      end
      12'b011010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1710;
      end
      12'b011010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1711;
      end
      12'b011010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1712;
      end
      12'b011010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1713;
      end
      12'b011010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1714;
      end
      12'b011010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1715;
      end
      12'b011010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1716;
      end
      12'b011010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1717;
      end
      12'b011010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1718;
      end
      12'b011010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1719;
      end
      12'b011010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1720;
      end
      12'b011010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1721;
      end
      12'b011010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1722;
      end
      12'b011010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1723;
      end
      12'b011010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1724;
      end
      12'b011010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1725;
      end
      12'b011010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1726;
      end
      12'b011010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1727;
      end
      12'b011011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1728;
      end
      12'b011011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1729;
      end
      12'b011011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1730;
      end
      12'b011011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1731;
      end
      12'b011011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1732;
      end
      12'b011011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1733;
      end
      12'b011011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1734;
      end
      12'b011011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1735;
      end
      12'b011011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1736;
      end
      12'b011011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1737;
      end
      12'b011011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1738;
      end
      12'b011011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1739;
      end
      12'b011011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1740;
      end
      12'b011011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1741;
      end
      12'b011011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1742;
      end
      12'b011011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1743;
      end
      12'b011011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1744;
      end
      12'b011011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1745;
      end
      12'b011011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1746;
      end
      12'b011011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1747;
      end
      12'b011011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1748;
      end
      12'b011011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1749;
      end
      12'b011011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1750;
      end
      12'b011011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1751;
      end
      12'b011011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1752;
      end
      12'b011011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1753;
      end
      12'b011011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1754;
      end
      12'b011011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1755;
      end
      12'b011011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1756;
      end
      12'b011011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1757;
      end
      12'b011011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1758;
      end
      12'b011011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1759;
      end
      12'b011011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1760;
      end
      12'b011011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1761;
      end
      12'b011011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1762;
      end
      12'b011011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1763;
      end
      12'b011011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1764;
      end
      12'b011011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1765;
      end
      12'b011011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1766;
      end
      12'b011011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1767;
      end
      12'b011011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1768;
      end
      12'b011011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1769;
      end
      12'b011011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1770;
      end
      12'b011011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1771;
      end
      12'b011011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1772;
      end
      12'b011011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1773;
      end
      12'b011011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1774;
      end
      12'b011011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1775;
      end
      12'b011011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1776;
      end
      12'b011011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1777;
      end
      12'b011011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1778;
      end
      12'b011011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1779;
      end
      12'b011011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1780;
      end
      12'b011011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1781;
      end
      12'b011011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1782;
      end
      12'b011011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1783;
      end
      12'b011011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1784;
      end
      12'b011011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1785;
      end
      12'b011011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1786;
      end
      12'b011011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1787;
      end
      12'b011011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1788;
      end
      12'b011011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1789;
      end
      12'b011011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1790;
      end
      12'b011011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1791;
      end
      12'b011100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1792;
      end
      12'b011100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1793;
      end
      12'b011100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1794;
      end
      12'b011100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1795;
      end
      12'b011100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1796;
      end
      12'b011100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1797;
      end
      12'b011100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1798;
      end
      12'b011100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1799;
      end
      12'b011100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1800;
      end
      12'b011100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1801;
      end
      12'b011100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1802;
      end
      12'b011100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1803;
      end
      12'b011100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1804;
      end
      12'b011100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1805;
      end
      12'b011100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1806;
      end
      12'b011100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1807;
      end
      12'b011100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1808;
      end
      12'b011100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1809;
      end
      12'b011100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1810;
      end
      12'b011100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1811;
      end
      12'b011100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1812;
      end
      12'b011100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1813;
      end
      12'b011100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1814;
      end
      12'b011100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1815;
      end
      12'b011100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1816;
      end
      12'b011100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1817;
      end
      12'b011100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1818;
      end
      12'b011100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1819;
      end
      12'b011100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1820;
      end
      12'b011100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1821;
      end
      12'b011100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1822;
      end
      12'b011100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1823;
      end
      12'b011100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1824;
      end
      12'b011100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1825;
      end
      12'b011100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1826;
      end
      12'b011100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1827;
      end
      12'b011100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1828;
      end
      12'b011100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1829;
      end
      12'b011100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1830;
      end
      12'b011100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1831;
      end
      12'b011100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1832;
      end
      12'b011100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1833;
      end
      12'b011100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1834;
      end
      12'b011100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1835;
      end
      12'b011100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1836;
      end
      12'b011100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1837;
      end
      12'b011100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1838;
      end
      12'b011100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1839;
      end
      12'b011100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1840;
      end
      12'b011100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1841;
      end
      12'b011100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1842;
      end
      12'b011100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1843;
      end
      12'b011100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1844;
      end
      12'b011100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1845;
      end
      12'b011100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1846;
      end
      12'b011100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1847;
      end
      12'b011100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1848;
      end
      12'b011100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1849;
      end
      12'b011100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1850;
      end
      12'b011100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1851;
      end
      12'b011100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1852;
      end
      12'b011100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1853;
      end
      12'b011100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1854;
      end
      12'b011100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1855;
      end
      12'b011101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1856;
      end
      12'b011101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1857;
      end
      12'b011101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1858;
      end
      12'b011101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1859;
      end
      12'b011101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1860;
      end
      12'b011101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1861;
      end
      12'b011101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1862;
      end
      12'b011101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1863;
      end
      12'b011101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1864;
      end
      12'b011101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1865;
      end
      12'b011101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1866;
      end
      12'b011101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1867;
      end
      12'b011101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1868;
      end
      12'b011101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1869;
      end
      12'b011101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1870;
      end
      12'b011101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1871;
      end
      12'b011101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1872;
      end
      12'b011101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1873;
      end
      12'b011101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1874;
      end
      12'b011101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1875;
      end
      12'b011101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1876;
      end
      12'b011101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1877;
      end
      12'b011101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1878;
      end
      12'b011101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1879;
      end
      12'b011101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1880;
      end
      12'b011101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1881;
      end
      12'b011101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1882;
      end
      12'b011101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1883;
      end
      12'b011101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1884;
      end
      12'b011101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1885;
      end
      12'b011101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1886;
      end
      12'b011101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1887;
      end
      12'b011101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1888;
      end
      12'b011101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1889;
      end
      12'b011101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1890;
      end
      12'b011101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1891;
      end
      12'b011101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1892;
      end
      12'b011101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1893;
      end
      12'b011101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1894;
      end
      12'b011101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1895;
      end
      12'b011101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1896;
      end
      12'b011101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1897;
      end
      12'b011101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1898;
      end
      12'b011101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1899;
      end
      12'b011101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1900;
      end
      12'b011101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1901;
      end
      12'b011101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1902;
      end
      12'b011101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1903;
      end
      12'b011101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1904;
      end
      12'b011101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1905;
      end
      12'b011101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1906;
      end
      12'b011101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1907;
      end
      12'b011101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1908;
      end
      12'b011101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1909;
      end
      12'b011101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1910;
      end
      12'b011101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1911;
      end
      12'b011101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1912;
      end
      12'b011101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1913;
      end
      12'b011101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1914;
      end
      12'b011101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1915;
      end
      12'b011101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1916;
      end
      12'b011101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1917;
      end
      12'b011101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1918;
      end
      12'b011101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1919;
      end
      12'b011110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1920;
      end
      12'b011110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1921;
      end
      12'b011110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1922;
      end
      12'b011110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1923;
      end
      12'b011110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1924;
      end
      12'b011110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1925;
      end
      12'b011110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1926;
      end
      12'b011110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1927;
      end
      12'b011110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1928;
      end
      12'b011110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1929;
      end
      12'b011110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1930;
      end
      12'b011110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1931;
      end
      12'b011110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1932;
      end
      12'b011110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1933;
      end
      12'b011110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1934;
      end
      12'b011110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1935;
      end
      12'b011110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_1936;
      end
      12'b011110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_1937;
      end
      12'b011110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_1938;
      end
      12'b011110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_1939;
      end
      12'b011110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_1940;
      end
      12'b011110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_1941;
      end
      12'b011110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_1942;
      end
      12'b011110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_1943;
      end
      12'b011110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_1944;
      end
      12'b011110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_1945;
      end
      12'b011110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_1946;
      end
      12'b011110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_1947;
      end
      12'b011110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_1948;
      end
      12'b011110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_1949;
      end
      12'b011110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_1950;
      end
      12'b011110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_1951;
      end
      12'b011110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_1952;
      end
      12'b011110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_1953;
      end
      12'b011110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_1954;
      end
      12'b011110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_1955;
      end
      12'b011110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_1956;
      end
      12'b011110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_1957;
      end
      12'b011110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_1958;
      end
      12'b011110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_1959;
      end
      12'b011110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_1960;
      end
      12'b011110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_1961;
      end
      12'b011110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_1962;
      end
      12'b011110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_1963;
      end
      12'b011110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_1964;
      end
      12'b011110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_1965;
      end
      12'b011110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_1966;
      end
      12'b011110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_1967;
      end
      12'b011110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_1968;
      end
      12'b011110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_1969;
      end
      12'b011110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_1970;
      end
      12'b011110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_1971;
      end
      12'b011110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_1972;
      end
      12'b011110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_1973;
      end
      12'b011110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_1974;
      end
      12'b011110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_1975;
      end
      12'b011110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_1976;
      end
      12'b011110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_1977;
      end
      12'b011110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_1978;
      end
      12'b011110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_1979;
      end
      12'b011110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_1980;
      end
      12'b011110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_1981;
      end
      12'b011110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_1982;
      end
      12'b011110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_1983;
      end
      12'b011111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_1984;
      end
      12'b011111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_1985;
      end
      12'b011111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_1986;
      end
      12'b011111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_1987;
      end
      12'b011111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_1988;
      end
      12'b011111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_1989;
      end
      12'b011111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_1990;
      end
      12'b011111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_1991;
      end
      12'b011111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_1992;
      end
      12'b011111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_1993;
      end
      12'b011111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_1994;
      end
      12'b011111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_1995;
      end
      12'b011111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_1996;
      end
      12'b011111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_1997;
      end
      12'b011111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_1998;
      end
      12'b011111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_1999;
      end
      12'b011111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2000;
      end
      12'b011111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2001;
      end
      12'b011111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2002;
      end
      12'b011111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2003;
      end
      12'b011111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2004;
      end
      12'b011111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2005;
      end
      12'b011111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2006;
      end
      12'b011111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2007;
      end
      12'b011111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2008;
      end
      12'b011111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2009;
      end
      12'b011111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2010;
      end
      12'b011111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2011;
      end
      12'b011111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2012;
      end
      12'b011111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2013;
      end
      12'b011111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2014;
      end
      12'b011111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2015;
      end
      12'b011111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2016;
      end
      12'b011111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2017;
      end
      12'b011111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2018;
      end
      12'b011111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2019;
      end
      12'b011111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2020;
      end
      12'b011111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2021;
      end
      12'b011111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2022;
      end
      12'b011111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2023;
      end
      12'b011111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2024;
      end
      12'b011111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2025;
      end
      12'b011111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2026;
      end
      12'b011111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2027;
      end
      12'b011111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2028;
      end
      12'b011111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2029;
      end
      12'b011111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2030;
      end
      12'b011111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2031;
      end
      12'b011111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2032;
      end
      12'b011111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2033;
      end
      12'b011111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2034;
      end
      12'b011111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2035;
      end
      12'b011111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2036;
      end
      12'b011111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2037;
      end
      12'b011111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2038;
      end
      12'b011111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2039;
      end
      12'b011111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2040;
      end
      12'b011111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2041;
      end
      12'b011111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2042;
      end
      12'b011111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2043;
      end
      12'b011111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2044;
      end
      12'b011111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2045;
      end
      12'b011111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2046;
      end
      12'b011111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2047;
      end
      12'b100000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2048;
      end
      12'b100000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2049;
      end
      12'b100000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2050;
      end
      12'b100000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2051;
      end
      12'b100000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2052;
      end
      12'b100000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2053;
      end
      12'b100000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2054;
      end
      12'b100000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2055;
      end
      12'b100000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2056;
      end
      12'b100000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2057;
      end
      12'b100000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2058;
      end
      12'b100000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2059;
      end
      12'b100000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2060;
      end
      12'b100000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2061;
      end
      12'b100000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2062;
      end
      12'b100000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2063;
      end
      12'b100000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2064;
      end
      12'b100000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2065;
      end
      12'b100000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2066;
      end
      12'b100000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2067;
      end
      12'b100000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2068;
      end
      12'b100000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2069;
      end
      12'b100000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2070;
      end
      12'b100000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2071;
      end
      12'b100000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2072;
      end
      12'b100000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2073;
      end
      12'b100000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2074;
      end
      12'b100000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2075;
      end
      12'b100000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2076;
      end
      12'b100000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2077;
      end
      12'b100000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2078;
      end
      12'b100000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2079;
      end
      12'b100000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2080;
      end
      12'b100000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2081;
      end
      12'b100000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2082;
      end
      12'b100000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2083;
      end
      12'b100000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2084;
      end
      12'b100000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2085;
      end
      12'b100000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2086;
      end
      12'b100000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2087;
      end
      12'b100000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2088;
      end
      12'b100000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2089;
      end
      12'b100000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2090;
      end
      12'b100000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2091;
      end
      12'b100000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2092;
      end
      12'b100000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2093;
      end
      12'b100000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2094;
      end
      12'b100000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2095;
      end
      12'b100000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2096;
      end
      12'b100000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2097;
      end
      12'b100000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2098;
      end
      12'b100000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2099;
      end
      12'b100000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2100;
      end
      12'b100000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2101;
      end
      12'b100000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2102;
      end
      12'b100000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2103;
      end
      12'b100000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2104;
      end
      12'b100000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2105;
      end
      12'b100000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2106;
      end
      12'b100000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2107;
      end
      12'b100000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2108;
      end
      12'b100000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2109;
      end
      12'b100000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2110;
      end
      12'b100000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2111;
      end
      12'b100001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2112;
      end
      12'b100001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2113;
      end
      12'b100001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2114;
      end
      12'b100001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2115;
      end
      12'b100001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2116;
      end
      12'b100001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2117;
      end
      12'b100001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2118;
      end
      12'b100001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2119;
      end
      12'b100001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2120;
      end
      12'b100001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2121;
      end
      12'b100001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2122;
      end
      12'b100001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2123;
      end
      12'b100001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2124;
      end
      12'b100001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2125;
      end
      12'b100001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2126;
      end
      12'b100001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2127;
      end
      12'b100001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2128;
      end
      12'b100001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2129;
      end
      12'b100001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2130;
      end
      12'b100001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2131;
      end
      12'b100001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2132;
      end
      12'b100001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2133;
      end
      12'b100001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2134;
      end
      12'b100001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2135;
      end
      12'b100001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2136;
      end
      12'b100001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2137;
      end
      12'b100001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2138;
      end
      12'b100001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2139;
      end
      12'b100001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2140;
      end
      12'b100001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2141;
      end
      12'b100001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2142;
      end
      12'b100001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2143;
      end
      12'b100001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2144;
      end
      12'b100001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2145;
      end
      12'b100001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2146;
      end
      12'b100001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2147;
      end
      12'b100001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2148;
      end
      12'b100001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2149;
      end
      12'b100001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2150;
      end
      12'b100001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2151;
      end
      12'b100001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2152;
      end
      12'b100001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2153;
      end
      12'b100001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2154;
      end
      12'b100001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2155;
      end
      12'b100001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2156;
      end
      12'b100001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2157;
      end
      12'b100001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2158;
      end
      12'b100001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2159;
      end
      12'b100001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2160;
      end
      12'b100001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2161;
      end
      12'b100001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2162;
      end
      12'b100001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2163;
      end
      12'b100001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2164;
      end
      12'b100001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2165;
      end
      12'b100001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2166;
      end
      12'b100001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2167;
      end
      12'b100001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2168;
      end
      12'b100001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2169;
      end
      12'b100001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2170;
      end
      12'b100001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2171;
      end
      12'b100001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2172;
      end
      12'b100001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2173;
      end
      12'b100001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2174;
      end
      12'b100001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2175;
      end
      12'b100010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2176;
      end
      12'b100010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2177;
      end
      12'b100010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2178;
      end
      12'b100010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2179;
      end
      12'b100010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2180;
      end
      12'b100010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2181;
      end
      12'b100010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2182;
      end
      12'b100010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2183;
      end
      12'b100010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2184;
      end
      12'b100010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2185;
      end
      12'b100010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2186;
      end
      12'b100010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2187;
      end
      12'b100010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2188;
      end
      12'b100010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2189;
      end
      12'b100010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2190;
      end
      12'b100010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2191;
      end
      12'b100010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2192;
      end
      12'b100010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2193;
      end
      12'b100010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2194;
      end
      12'b100010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2195;
      end
      12'b100010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2196;
      end
      12'b100010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2197;
      end
      12'b100010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2198;
      end
      12'b100010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2199;
      end
      12'b100010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2200;
      end
      12'b100010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2201;
      end
      12'b100010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2202;
      end
      12'b100010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2203;
      end
      12'b100010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2204;
      end
      12'b100010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2205;
      end
      12'b100010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2206;
      end
      12'b100010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2207;
      end
      12'b100010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2208;
      end
      12'b100010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2209;
      end
      12'b100010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2210;
      end
      12'b100010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2211;
      end
      12'b100010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2212;
      end
      12'b100010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2213;
      end
      12'b100010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2214;
      end
      12'b100010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2215;
      end
      12'b100010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2216;
      end
      12'b100010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2217;
      end
      12'b100010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2218;
      end
      12'b100010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2219;
      end
      12'b100010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2220;
      end
      12'b100010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2221;
      end
      12'b100010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2222;
      end
      12'b100010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2223;
      end
      12'b100010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2224;
      end
      12'b100010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2225;
      end
      12'b100010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2226;
      end
      12'b100010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2227;
      end
      12'b100010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2228;
      end
      12'b100010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2229;
      end
      12'b100010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2230;
      end
      12'b100010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2231;
      end
      12'b100010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2232;
      end
      12'b100010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2233;
      end
      12'b100010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2234;
      end
      12'b100010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2235;
      end
      12'b100010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2236;
      end
      12'b100010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2237;
      end
      12'b100010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2238;
      end
      12'b100010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2239;
      end
      12'b100011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2240;
      end
      12'b100011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2241;
      end
      12'b100011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2242;
      end
      12'b100011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2243;
      end
      12'b100011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2244;
      end
      12'b100011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2245;
      end
      12'b100011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2246;
      end
      12'b100011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2247;
      end
      12'b100011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2248;
      end
      12'b100011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2249;
      end
      12'b100011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2250;
      end
      12'b100011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2251;
      end
      12'b100011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2252;
      end
      12'b100011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2253;
      end
      12'b100011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2254;
      end
      12'b100011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2255;
      end
      12'b100011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2256;
      end
      12'b100011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2257;
      end
      12'b100011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2258;
      end
      12'b100011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2259;
      end
      12'b100011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2260;
      end
      12'b100011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2261;
      end
      12'b100011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2262;
      end
      12'b100011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2263;
      end
      12'b100011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2264;
      end
      12'b100011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2265;
      end
      12'b100011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2266;
      end
      12'b100011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2267;
      end
      12'b100011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2268;
      end
      12'b100011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2269;
      end
      12'b100011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2270;
      end
      12'b100011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2271;
      end
      12'b100011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2272;
      end
      12'b100011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2273;
      end
      12'b100011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2274;
      end
      12'b100011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2275;
      end
      12'b100011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2276;
      end
      12'b100011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2277;
      end
      12'b100011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2278;
      end
      12'b100011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2279;
      end
      12'b100011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2280;
      end
      12'b100011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2281;
      end
      12'b100011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2282;
      end
      12'b100011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2283;
      end
      12'b100011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2284;
      end
      12'b100011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2285;
      end
      12'b100011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2286;
      end
      12'b100011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2287;
      end
      12'b100011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2288;
      end
      12'b100011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2289;
      end
      12'b100011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2290;
      end
      12'b100011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2291;
      end
      12'b100011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2292;
      end
      12'b100011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2293;
      end
      12'b100011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2294;
      end
      12'b100011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2295;
      end
      12'b100011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2296;
      end
      12'b100011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2297;
      end
      12'b100011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2298;
      end
      12'b100011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2299;
      end
      12'b100011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2300;
      end
      12'b100011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2301;
      end
      12'b100011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2302;
      end
      12'b100011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2303;
      end
      12'b100100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2304;
      end
      12'b100100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2305;
      end
      12'b100100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2306;
      end
      12'b100100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2307;
      end
      12'b100100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2308;
      end
      12'b100100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2309;
      end
      12'b100100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2310;
      end
      12'b100100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2311;
      end
      12'b100100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2312;
      end
      12'b100100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2313;
      end
      12'b100100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2314;
      end
      12'b100100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2315;
      end
      12'b100100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2316;
      end
      12'b100100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2317;
      end
      12'b100100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2318;
      end
      12'b100100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2319;
      end
      12'b100100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2320;
      end
      12'b100100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2321;
      end
      12'b100100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2322;
      end
      12'b100100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2323;
      end
      12'b100100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2324;
      end
      12'b100100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2325;
      end
      12'b100100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2326;
      end
      12'b100100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2327;
      end
      12'b100100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2328;
      end
      12'b100100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2329;
      end
      12'b100100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2330;
      end
      12'b100100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2331;
      end
      12'b100100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2332;
      end
      12'b100100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2333;
      end
      12'b100100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2334;
      end
      12'b100100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2335;
      end
      12'b100100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2336;
      end
      12'b100100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2337;
      end
      12'b100100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2338;
      end
      12'b100100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2339;
      end
      12'b100100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2340;
      end
      12'b100100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2341;
      end
      12'b100100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2342;
      end
      12'b100100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2343;
      end
      12'b100100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2344;
      end
      12'b100100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2345;
      end
      12'b100100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2346;
      end
      12'b100100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2347;
      end
      12'b100100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2348;
      end
      12'b100100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2349;
      end
      12'b100100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2350;
      end
      12'b100100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2351;
      end
      12'b100100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2352;
      end
      12'b100100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2353;
      end
      12'b100100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2354;
      end
      12'b100100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2355;
      end
      12'b100100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2356;
      end
      12'b100100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2357;
      end
      12'b100100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2358;
      end
      12'b100100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2359;
      end
      12'b100100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2360;
      end
      12'b100100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2361;
      end
      12'b100100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2362;
      end
      12'b100100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2363;
      end
      12'b100100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2364;
      end
      12'b100100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2365;
      end
      12'b100100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2366;
      end
      12'b100100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2367;
      end
      12'b100101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2368;
      end
      12'b100101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2369;
      end
      12'b100101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2370;
      end
      12'b100101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2371;
      end
      12'b100101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2372;
      end
      12'b100101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2373;
      end
      12'b100101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2374;
      end
      12'b100101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2375;
      end
      12'b100101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2376;
      end
      12'b100101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2377;
      end
      12'b100101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2378;
      end
      12'b100101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2379;
      end
      12'b100101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2380;
      end
      12'b100101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2381;
      end
      12'b100101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2382;
      end
      12'b100101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2383;
      end
      12'b100101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2384;
      end
      12'b100101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2385;
      end
      12'b100101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2386;
      end
      12'b100101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2387;
      end
      12'b100101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2388;
      end
      12'b100101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2389;
      end
      12'b100101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2390;
      end
      12'b100101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2391;
      end
      12'b100101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2392;
      end
      12'b100101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2393;
      end
      12'b100101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2394;
      end
      12'b100101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2395;
      end
      12'b100101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2396;
      end
      12'b100101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2397;
      end
      12'b100101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2398;
      end
      12'b100101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2399;
      end
      12'b100101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2400;
      end
      12'b100101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2401;
      end
      12'b100101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2402;
      end
      12'b100101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2403;
      end
      12'b100101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2404;
      end
      12'b100101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2405;
      end
      12'b100101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2406;
      end
      12'b100101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2407;
      end
      12'b100101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2408;
      end
      12'b100101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2409;
      end
      12'b100101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2410;
      end
      12'b100101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2411;
      end
      12'b100101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2412;
      end
      12'b100101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2413;
      end
      12'b100101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2414;
      end
      12'b100101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2415;
      end
      12'b100101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2416;
      end
      12'b100101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2417;
      end
      12'b100101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2418;
      end
      12'b100101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2419;
      end
      12'b100101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2420;
      end
      12'b100101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2421;
      end
      12'b100101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2422;
      end
      12'b100101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2423;
      end
      12'b100101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2424;
      end
      12'b100101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2425;
      end
      12'b100101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2426;
      end
      12'b100101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2427;
      end
      12'b100101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2428;
      end
      12'b100101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2429;
      end
      12'b100101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2430;
      end
      12'b100101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2431;
      end
      12'b100110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2432;
      end
      12'b100110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2433;
      end
      12'b100110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2434;
      end
      12'b100110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2435;
      end
      12'b100110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2436;
      end
      12'b100110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2437;
      end
      12'b100110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2438;
      end
      12'b100110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2439;
      end
      12'b100110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2440;
      end
      12'b100110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2441;
      end
      12'b100110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2442;
      end
      12'b100110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2443;
      end
      12'b100110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2444;
      end
      12'b100110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2445;
      end
      12'b100110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2446;
      end
      12'b100110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2447;
      end
      12'b100110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2448;
      end
      12'b100110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2449;
      end
      12'b100110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2450;
      end
      12'b100110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2451;
      end
      12'b100110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2452;
      end
      12'b100110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2453;
      end
      12'b100110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2454;
      end
      12'b100110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2455;
      end
      12'b100110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2456;
      end
      12'b100110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2457;
      end
      12'b100110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2458;
      end
      12'b100110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2459;
      end
      12'b100110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2460;
      end
      12'b100110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2461;
      end
      12'b100110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2462;
      end
      12'b100110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2463;
      end
      12'b100110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2464;
      end
      12'b100110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2465;
      end
      12'b100110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2466;
      end
      12'b100110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2467;
      end
      12'b100110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2468;
      end
      12'b100110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2469;
      end
      12'b100110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2470;
      end
      12'b100110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2471;
      end
      12'b100110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2472;
      end
      12'b100110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2473;
      end
      12'b100110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2474;
      end
      12'b100110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2475;
      end
      12'b100110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2476;
      end
      12'b100110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2477;
      end
      12'b100110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2478;
      end
      12'b100110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2479;
      end
      12'b100110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2480;
      end
      12'b100110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2481;
      end
      12'b100110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2482;
      end
      12'b100110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2483;
      end
      12'b100110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2484;
      end
      12'b100110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2485;
      end
      12'b100110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2486;
      end
      12'b100110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2487;
      end
      12'b100110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2488;
      end
      12'b100110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2489;
      end
      12'b100110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2490;
      end
      12'b100110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2491;
      end
      12'b100110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2492;
      end
      12'b100110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2493;
      end
      12'b100110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2494;
      end
      12'b100110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2495;
      end
      12'b100111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2496;
      end
      12'b100111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2497;
      end
      12'b100111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2498;
      end
      12'b100111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2499;
      end
      12'b100111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2500;
      end
      12'b100111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2501;
      end
      12'b100111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2502;
      end
      12'b100111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2503;
      end
      12'b100111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2504;
      end
      12'b100111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2505;
      end
      12'b100111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2506;
      end
      12'b100111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2507;
      end
      12'b100111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2508;
      end
      12'b100111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2509;
      end
      12'b100111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2510;
      end
      12'b100111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2511;
      end
      12'b100111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2512;
      end
      12'b100111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2513;
      end
      12'b100111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2514;
      end
      12'b100111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2515;
      end
      12'b100111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2516;
      end
      12'b100111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2517;
      end
      12'b100111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2518;
      end
      12'b100111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2519;
      end
      12'b100111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2520;
      end
      12'b100111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2521;
      end
      12'b100111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2522;
      end
      12'b100111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2523;
      end
      12'b100111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2524;
      end
      12'b100111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2525;
      end
      12'b100111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2526;
      end
      12'b100111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2527;
      end
      12'b100111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2528;
      end
      12'b100111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2529;
      end
      12'b100111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2530;
      end
      12'b100111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2531;
      end
      12'b100111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2532;
      end
      12'b100111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2533;
      end
      12'b100111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2534;
      end
      12'b100111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2535;
      end
      12'b100111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2536;
      end
      12'b100111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2537;
      end
      12'b100111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2538;
      end
      12'b100111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2539;
      end
      12'b100111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2540;
      end
      12'b100111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2541;
      end
      12'b100111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2542;
      end
      12'b100111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2543;
      end
      12'b100111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2544;
      end
      12'b100111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2545;
      end
      12'b100111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2546;
      end
      12'b100111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2547;
      end
      12'b100111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2548;
      end
      12'b100111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2549;
      end
      12'b100111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2550;
      end
      12'b100111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2551;
      end
      12'b100111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2552;
      end
      12'b100111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2553;
      end
      12'b100111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2554;
      end
      12'b100111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2555;
      end
      12'b100111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2556;
      end
      12'b100111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2557;
      end
      12'b100111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2558;
      end
      12'b100111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2559;
      end
      12'b101000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2560;
      end
      12'b101000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2561;
      end
      12'b101000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2562;
      end
      12'b101000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2563;
      end
      12'b101000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2564;
      end
      12'b101000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2565;
      end
      12'b101000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2566;
      end
      12'b101000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2567;
      end
      12'b101000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2568;
      end
      12'b101000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2569;
      end
      12'b101000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2570;
      end
      12'b101000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2571;
      end
      12'b101000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2572;
      end
      12'b101000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2573;
      end
      12'b101000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2574;
      end
      12'b101000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2575;
      end
      12'b101000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2576;
      end
      12'b101000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2577;
      end
      12'b101000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2578;
      end
      12'b101000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2579;
      end
      12'b101000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2580;
      end
      12'b101000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2581;
      end
      12'b101000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2582;
      end
      12'b101000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2583;
      end
      12'b101000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2584;
      end
      12'b101000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2585;
      end
      12'b101000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2586;
      end
      12'b101000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2587;
      end
      12'b101000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2588;
      end
      12'b101000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2589;
      end
      12'b101000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2590;
      end
      12'b101000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2591;
      end
      12'b101000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2592;
      end
      12'b101000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2593;
      end
      12'b101000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2594;
      end
      12'b101000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2595;
      end
      12'b101000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2596;
      end
      12'b101000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2597;
      end
      12'b101000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2598;
      end
      12'b101000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2599;
      end
      12'b101000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2600;
      end
      12'b101000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2601;
      end
      12'b101000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2602;
      end
      12'b101000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2603;
      end
      12'b101000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2604;
      end
      12'b101000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2605;
      end
      12'b101000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2606;
      end
      12'b101000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2607;
      end
      12'b101000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2608;
      end
      12'b101000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2609;
      end
      12'b101000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2610;
      end
      12'b101000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2611;
      end
      12'b101000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2612;
      end
      12'b101000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2613;
      end
      12'b101000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2614;
      end
      12'b101000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2615;
      end
      12'b101000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2616;
      end
      12'b101000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2617;
      end
      12'b101000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2618;
      end
      12'b101000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2619;
      end
      12'b101000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2620;
      end
      12'b101000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2621;
      end
      12'b101000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2622;
      end
      12'b101000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2623;
      end
      12'b101001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2624;
      end
      12'b101001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2625;
      end
      12'b101001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2626;
      end
      12'b101001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2627;
      end
      12'b101001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2628;
      end
      12'b101001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2629;
      end
      12'b101001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2630;
      end
      12'b101001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2631;
      end
      12'b101001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2632;
      end
      12'b101001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2633;
      end
      12'b101001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2634;
      end
      12'b101001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2635;
      end
      12'b101001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2636;
      end
      12'b101001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2637;
      end
      12'b101001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2638;
      end
      12'b101001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2639;
      end
      12'b101001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2640;
      end
      12'b101001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2641;
      end
      12'b101001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2642;
      end
      12'b101001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2643;
      end
      12'b101001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2644;
      end
      12'b101001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2645;
      end
      12'b101001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2646;
      end
      12'b101001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2647;
      end
      12'b101001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2648;
      end
      12'b101001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2649;
      end
      12'b101001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2650;
      end
      12'b101001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2651;
      end
      12'b101001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2652;
      end
      12'b101001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2653;
      end
      12'b101001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2654;
      end
      12'b101001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2655;
      end
      12'b101001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2656;
      end
      12'b101001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2657;
      end
      12'b101001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2658;
      end
      12'b101001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2659;
      end
      12'b101001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2660;
      end
      12'b101001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2661;
      end
      12'b101001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2662;
      end
      12'b101001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2663;
      end
      12'b101001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2664;
      end
      12'b101001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2665;
      end
      12'b101001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2666;
      end
      12'b101001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2667;
      end
      12'b101001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2668;
      end
      12'b101001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2669;
      end
      12'b101001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2670;
      end
      12'b101001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2671;
      end
      12'b101001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2672;
      end
      12'b101001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2673;
      end
      12'b101001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2674;
      end
      12'b101001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2675;
      end
      12'b101001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2676;
      end
      12'b101001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2677;
      end
      12'b101001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2678;
      end
      12'b101001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2679;
      end
      12'b101001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2680;
      end
      12'b101001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2681;
      end
      12'b101001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2682;
      end
      12'b101001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2683;
      end
      12'b101001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2684;
      end
      12'b101001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2685;
      end
      12'b101001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2686;
      end
      12'b101001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2687;
      end
      12'b101010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2688;
      end
      12'b101010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2689;
      end
      12'b101010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2690;
      end
      12'b101010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2691;
      end
      12'b101010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2692;
      end
      12'b101010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2693;
      end
      12'b101010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2694;
      end
      12'b101010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2695;
      end
      12'b101010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2696;
      end
      12'b101010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2697;
      end
      12'b101010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2698;
      end
      12'b101010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2699;
      end
      12'b101010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2700;
      end
      12'b101010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2701;
      end
      12'b101010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2702;
      end
      12'b101010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2703;
      end
      12'b101010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2704;
      end
      12'b101010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2705;
      end
      12'b101010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2706;
      end
      12'b101010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2707;
      end
      12'b101010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2708;
      end
      12'b101010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2709;
      end
      12'b101010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2710;
      end
      12'b101010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2711;
      end
      12'b101010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2712;
      end
      12'b101010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2713;
      end
      12'b101010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2714;
      end
      12'b101010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2715;
      end
      12'b101010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2716;
      end
      12'b101010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2717;
      end
      12'b101010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2718;
      end
      12'b101010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2719;
      end
      12'b101010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2720;
      end
      12'b101010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2721;
      end
      12'b101010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2722;
      end
      12'b101010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2723;
      end
      12'b101010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2724;
      end
      12'b101010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2725;
      end
      12'b101010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2726;
      end
      12'b101010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2727;
      end
      12'b101010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2728;
      end
      12'b101010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2729;
      end
      12'b101010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2730;
      end
      12'b101010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2731;
      end
      12'b101010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2732;
      end
      12'b101010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2733;
      end
      12'b101010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2734;
      end
      12'b101010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2735;
      end
      12'b101010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2736;
      end
      12'b101010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2737;
      end
      12'b101010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2738;
      end
      12'b101010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2739;
      end
      12'b101010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2740;
      end
      12'b101010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2741;
      end
      12'b101010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2742;
      end
      12'b101010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2743;
      end
      12'b101010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2744;
      end
      12'b101010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2745;
      end
      12'b101010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2746;
      end
      12'b101010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2747;
      end
      12'b101010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2748;
      end
      12'b101010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2749;
      end
      12'b101010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2750;
      end
      12'b101010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2751;
      end
      12'b101011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2752;
      end
      12'b101011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2753;
      end
      12'b101011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2754;
      end
      12'b101011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2755;
      end
      12'b101011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2756;
      end
      12'b101011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2757;
      end
      12'b101011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2758;
      end
      12'b101011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2759;
      end
      12'b101011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2760;
      end
      12'b101011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2761;
      end
      12'b101011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2762;
      end
      12'b101011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2763;
      end
      12'b101011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2764;
      end
      12'b101011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2765;
      end
      12'b101011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2766;
      end
      12'b101011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2767;
      end
      12'b101011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2768;
      end
      12'b101011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2769;
      end
      12'b101011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2770;
      end
      12'b101011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2771;
      end
      12'b101011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2772;
      end
      12'b101011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2773;
      end
      12'b101011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2774;
      end
      12'b101011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2775;
      end
      12'b101011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2776;
      end
      12'b101011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2777;
      end
      12'b101011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2778;
      end
      12'b101011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2779;
      end
      12'b101011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2780;
      end
      12'b101011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2781;
      end
      12'b101011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2782;
      end
      12'b101011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2783;
      end
      12'b101011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2784;
      end
      12'b101011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2785;
      end
      12'b101011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2786;
      end
      12'b101011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2787;
      end
      12'b101011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2788;
      end
      12'b101011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2789;
      end
      12'b101011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2790;
      end
      12'b101011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2791;
      end
      12'b101011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2792;
      end
      12'b101011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2793;
      end
      12'b101011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2794;
      end
      12'b101011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2795;
      end
      12'b101011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2796;
      end
      12'b101011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2797;
      end
      12'b101011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2798;
      end
      12'b101011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2799;
      end
      12'b101011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2800;
      end
      12'b101011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2801;
      end
      12'b101011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2802;
      end
      12'b101011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2803;
      end
      12'b101011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2804;
      end
      12'b101011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2805;
      end
      12'b101011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2806;
      end
      12'b101011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2807;
      end
      12'b101011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2808;
      end
      12'b101011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2809;
      end
      12'b101011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2810;
      end
      12'b101011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2811;
      end
      12'b101011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2812;
      end
      12'b101011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2813;
      end
      12'b101011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2814;
      end
      12'b101011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2815;
      end
      12'b101100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2816;
      end
      12'b101100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2817;
      end
      12'b101100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2818;
      end
      12'b101100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2819;
      end
      12'b101100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2820;
      end
      12'b101100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2821;
      end
      12'b101100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2822;
      end
      12'b101100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2823;
      end
      12'b101100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2824;
      end
      12'b101100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2825;
      end
      12'b101100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2826;
      end
      12'b101100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2827;
      end
      12'b101100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2828;
      end
      12'b101100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2829;
      end
      12'b101100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2830;
      end
      12'b101100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2831;
      end
      12'b101100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2832;
      end
      12'b101100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2833;
      end
      12'b101100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2834;
      end
      12'b101100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2835;
      end
      12'b101100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2836;
      end
      12'b101100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2837;
      end
      12'b101100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2838;
      end
      12'b101100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2839;
      end
      12'b101100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2840;
      end
      12'b101100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2841;
      end
      12'b101100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2842;
      end
      12'b101100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2843;
      end
      12'b101100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2844;
      end
      12'b101100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2845;
      end
      12'b101100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2846;
      end
      12'b101100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2847;
      end
      12'b101100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2848;
      end
      12'b101100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2849;
      end
      12'b101100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2850;
      end
      12'b101100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2851;
      end
      12'b101100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2852;
      end
      12'b101100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2853;
      end
      12'b101100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2854;
      end
      12'b101100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2855;
      end
      12'b101100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2856;
      end
      12'b101100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2857;
      end
      12'b101100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2858;
      end
      12'b101100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2859;
      end
      12'b101100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2860;
      end
      12'b101100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2861;
      end
      12'b101100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2862;
      end
      12'b101100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2863;
      end
      12'b101100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2864;
      end
      12'b101100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2865;
      end
      12'b101100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2866;
      end
      12'b101100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2867;
      end
      12'b101100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2868;
      end
      12'b101100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2869;
      end
      12'b101100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2870;
      end
      12'b101100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2871;
      end
      12'b101100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2872;
      end
      12'b101100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2873;
      end
      12'b101100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2874;
      end
      12'b101100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2875;
      end
      12'b101100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2876;
      end
      12'b101100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2877;
      end
      12'b101100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2878;
      end
      12'b101100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2879;
      end
      12'b101101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2880;
      end
      12'b101101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2881;
      end
      12'b101101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2882;
      end
      12'b101101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2883;
      end
      12'b101101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2884;
      end
      12'b101101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2885;
      end
      12'b101101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2886;
      end
      12'b101101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2887;
      end
      12'b101101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2888;
      end
      12'b101101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2889;
      end
      12'b101101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2890;
      end
      12'b101101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2891;
      end
      12'b101101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2892;
      end
      12'b101101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2893;
      end
      12'b101101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2894;
      end
      12'b101101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2895;
      end
      12'b101101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2896;
      end
      12'b101101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2897;
      end
      12'b101101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2898;
      end
      12'b101101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2899;
      end
      12'b101101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2900;
      end
      12'b101101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2901;
      end
      12'b101101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2902;
      end
      12'b101101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2903;
      end
      12'b101101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2904;
      end
      12'b101101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2905;
      end
      12'b101101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2906;
      end
      12'b101101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2907;
      end
      12'b101101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2908;
      end
      12'b101101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2909;
      end
      12'b101101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2910;
      end
      12'b101101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2911;
      end
      12'b101101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2912;
      end
      12'b101101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2913;
      end
      12'b101101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2914;
      end
      12'b101101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2915;
      end
      12'b101101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2916;
      end
      12'b101101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2917;
      end
      12'b101101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2918;
      end
      12'b101101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2919;
      end
      12'b101101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2920;
      end
      12'b101101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2921;
      end
      12'b101101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2922;
      end
      12'b101101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2923;
      end
      12'b101101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2924;
      end
      12'b101101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2925;
      end
      12'b101101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2926;
      end
      12'b101101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2927;
      end
      12'b101101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2928;
      end
      12'b101101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2929;
      end
      12'b101101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2930;
      end
      12'b101101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2931;
      end
      12'b101101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2932;
      end
      12'b101101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2933;
      end
      12'b101101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2934;
      end
      12'b101101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2935;
      end
      12'b101101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_2936;
      end
      12'b101101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_2937;
      end
      12'b101101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_2938;
      end
      12'b101101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_2939;
      end
      12'b101101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_2940;
      end
      12'b101101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_2941;
      end
      12'b101101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_2942;
      end
      12'b101101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_2943;
      end
      12'b101110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_2944;
      end
      12'b101110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_2945;
      end
      12'b101110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_2946;
      end
      12'b101110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_2947;
      end
      12'b101110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_2948;
      end
      12'b101110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_2949;
      end
      12'b101110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_2950;
      end
      12'b101110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_2951;
      end
      12'b101110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_2952;
      end
      12'b101110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_2953;
      end
      12'b101110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_2954;
      end
      12'b101110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_2955;
      end
      12'b101110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_2956;
      end
      12'b101110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_2957;
      end
      12'b101110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_2958;
      end
      12'b101110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_2959;
      end
      12'b101110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_2960;
      end
      12'b101110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_2961;
      end
      12'b101110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_2962;
      end
      12'b101110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_2963;
      end
      12'b101110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_2964;
      end
      12'b101110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_2965;
      end
      12'b101110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_2966;
      end
      12'b101110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_2967;
      end
      12'b101110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_2968;
      end
      12'b101110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_2969;
      end
      12'b101110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_2970;
      end
      12'b101110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_2971;
      end
      12'b101110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_2972;
      end
      12'b101110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_2973;
      end
      12'b101110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_2974;
      end
      12'b101110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_2975;
      end
      12'b101110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_2976;
      end
      12'b101110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_2977;
      end
      12'b101110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_2978;
      end
      12'b101110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_2979;
      end
      12'b101110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_2980;
      end
      12'b101110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_2981;
      end
      12'b101110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_2982;
      end
      12'b101110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_2983;
      end
      12'b101110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_2984;
      end
      12'b101110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_2985;
      end
      12'b101110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_2986;
      end
      12'b101110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_2987;
      end
      12'b101110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_2988;
      end
      12'b101110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_2989;
      end
      12'b101110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_2990;
      end
      12'b101110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_2991;
      end
      12'b101110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_2992;
      end
      12'b101110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_2993;
      end
      12'b101110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_2994;
      end
      12'b101110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_2995;
      end
      12'b101110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_2996;
      end
      12'b101110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_2997;
      end
      12'b101110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_2998;
      end
      12'b101110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_2999;
      end
      12'b101110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3000;
      end
      12'b101110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3001;
      end
      12'b101110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3002;
      end
      12'b101110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3003;
      end
      12'b101110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3004;
      end
      12'b101110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3005;
      end
      12'b101110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3006;
      end
      12'b101110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3007;
      end
      12'b101111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3008;
      end
      12'b101111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3009;
      end
      12'b101111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3010;
      end
      12'b101111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3011;
      end
      12'b101111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3012;
      end
      12'b101111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3013;
      end
      12'b101111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3014;
      end
      12'b101111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3015;
      end
      12'b101111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3016;
      end
      12'b101111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3017;
      end
      12'b101111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3018;
      end
      12'b101111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3019;
      end
      12'b101111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3020;
      end
      12'b101111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3021;
      end
      12'b101111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3022;
      end
      12'b101111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3023;
      end
      12'b101111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3024;
      end
      12'b101111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3025;
      end
      12'b101111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3026;
      end
      12'b101111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3027;
      end
      12'b101111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3028;
      end
      12'b101111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3029;
      end
      12'b101111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3030;
      end
      12'b101111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3031;
      end
      12'b101111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3032;
      end
      12'b101111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3033;
      end
      12'b101111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3034;
      end
      12'b101111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3035;
      end
      12'b101111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3036;
      end
      12'b101111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3037;
      end
      12'b101111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3038;
      end
      12'b101111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3039;
      end
      12'b101111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3040;
      end
      12'b101111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3041;
      end
      12'b101111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3042;
      end
      12'b101111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3043;
      end
      12'b101111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3044;
      end
      12'b101111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3045;
      end
      12'b101111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3046;
      end
      12'b101111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3047;
      end
      12'b101111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3048;
      end
      12'b101111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3049;
      end
      12'b101111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3050;
      end
      12'b101111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3051;
      end
      12'b101111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3052;
      end
      12'b101111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3053;
      end
      12'b101111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3054;
      end
      12'b101111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3055;
      end
      12'b101111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3056;
      end
      12'b101111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3057;
      end
      12'b101111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3058;
      end
      12'b101111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3059;
      end
      12'b101111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3060;
      end
      12'b101111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3061;
      end
      12'b101111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3062;
      end
      12'b101111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3063;
      end
      12'b101111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3064;
      end
      12'b101111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3065;
      end
      12'b101111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3066;
      end
      12'b101111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3067;
      end
      12'b101111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3068;
      end
      12'b101111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3069;
      end
      12'b101111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3070;
      end
      12'b101111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3071;
      end
      12'b110000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3072;
      end
      12'b110000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3073;
      end
      12'b110000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3074;
      end
      12'b110000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3075;
      end
      12'b110000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3076;
      end
      12'b110000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3077;
      end
      12'b110000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3078;
      end
      12'b110000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3079;
      end
      12'b110000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3080;
      end
      12'b110000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3081;
      end
      12'b110000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3082;
      end
      12'b110000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3083;
      end
      12'b110000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3084;
      end
      12'b110000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3085;
      end
      12'b110000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3086;
      end
      12'b110000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3087;
      end
      12'b110000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3088;
      end
      12'b110000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3089;
      end
      12'b110000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3090;
      end
      12'b110000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3091;
      end
      12'b110000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3092;
      end
      12'b110000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3093;
      end
      12'b110000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3094;
      end
      12'b110000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3095;
      end
      12'b110000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3096;
      end
      12'b110000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3097;
      end
      12'b110000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3098;
      end
      12'b110000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3099;
      end
      12'b110000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3100;
      end
      12'b110000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3101;
      end
      12'b110000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3102;
      end
      12'b110000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3103;
      end
      12'b110000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3104;
      end
      12'b110000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3105;
      end
      12'b110000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3106;
      end
      12'b110000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3107;
      end
      12'b110000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3108;
      end
      12'b110000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3109;
      end
      12'b110000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3110;
      end
      12'b110000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3111;
      end
      12'b110000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3112;
      end
      12'b110000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3113;
      end
      12'b110000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3114;
      end
      12'b110000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3115;
      end
      12'b110000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3116;
      end
      12'b110000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3117;
      end
      12'b110000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3118;
      end
      12'b110000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3119;
      end
      12'b110000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3120;
      end
      12'b110000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3121;
      end
      12'b110000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3122;
      end
      12'b110000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3123;
      end
      12'b110000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3124;
      end
      12'b110000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3125;
      end
      12'b110000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3126;
      end
      12'b110000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3127;
      end
      12'b110000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3128;
      end
      12'b110000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3129;
      end
      12'b110000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3130;
      end
      12'b110000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3131;
      end
      12'b110000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3132;
      end
      12'b110000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3133;
      end
      12'b110000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3134;
      end
      12'b110000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3135;
      end
      12'b110001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3136;
      end
      12'b110001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3137;
      end
      12'b110001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3138;
      end
      12'b110001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3139;
      end
      12'b110001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3140;
      end
      12'b110001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3141;
      end
      12'b110001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3142;
      end
      12'b110001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3143;
      end
      12'b110001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3144;
      end
      12'b110001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3145;
      end
      12'b110001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3146;
      end
      12'b110001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3147;
      end
      12'b110001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3148;
      end
      12'b110001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3149;
      end
      12'b110001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3150;
      end
      12'b110001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3151;
      end
      12'b110001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3152;
      end
      12'b110001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3153;
      end
      12'b110001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3154;
      end
      12'b110001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3155;
      end
      12'b110001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3156;
      end
      12'b110001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3157;
      end
      12'b110001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3158;
      end
      12'b110001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3159;
      end
      12'b110001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3160;
      end
      12'b110001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3161;
      end
      12'b110001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3162;
      end
      12'b110001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3163;
      end
      12'b110001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3164;
      end
      12'b110001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3165;
      end
      12'b110001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3166;
      end
      12'b110001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3167;
      end
      12'b110001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3168;
      end
      12'b110001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3169;
      end
      12'b110001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3170;
      end
      12'b110001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3171;
      end
      12'b110001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3172;
      end
      12'b110001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3173;
      end
      12'b110001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3174;
      end
      12'b110001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3175;
      end
      12'b110001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3176;
      end
      12'b110001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3177;
      end
      12'b110001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3178;
      end
      12'b110001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3179;
      end
      12'b110001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3180;
      end
      12'b110001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3181;
      end
      12'b110001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3182;
      end
      12'b110001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3183;
      end
      12'b110001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3184;
      end
      12'b110001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3185;
      end
      12'b110001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3186;
      end
      12'b110001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3187;
      end
      12'b110001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3188;
      end
      12'b110001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3189;
      end
      12'b110001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3190;
      end
      12'b110001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3191;
      end
      12'b110001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3192;
      end
      12'b110001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3193;
      end
      12'b110001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3194;
      end
      12'b110001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3195;
      end
      12'b110001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3196;
      end
      12'b110001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3197;
      end
      12'b110001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3198;
      end
      12'b110001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3199;
      end
      12'b110010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3200;
      end
      12'b110010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3201;
      end
      12'b110010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3202;
      end
      12'b110010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3203;
      end
      12'b110010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3204;
      end
      12'b110010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3205;
      end
      12'b110010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3206;
      end
      12'b110010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3207;
      end
      12'b110010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3208;
      end
      12'b110010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3209;
      end
      12'b110010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3210;
      end
      12'b110010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3211;
      end
      12'b110010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3212;
      end
      12'b110010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3213;
      end
      12'b110010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3214;
      end
      12'b110010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3215;
      end
      12'b110010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3216;
      end
      12'b110010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3217;
      end
      12'b110010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3218;
      end
      12'b110010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3219;
      end
      12'b110010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3220;
      end
      12'b110010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3221;
      end
      12'b110010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3222;
      end
      12'b110010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3223;
      end
      12'b110010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3224;
      end
      12'b110010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3225;
      end
      12'b110010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3226;
      end
      12'b110010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3227;
      end
      12'b110010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3228;
      end
      12'b110010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3229;
      end
      12'b110010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3230;
      end
      12'b110010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3231;
      end
      12'b110010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3232;
      end
      12'b110010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3233;
      end
      12'b110010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3234;
      end
      12'b110010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3235;
      end
      12'b110010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3236;
      end
      12'b110010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3237;
      end
      12'b110010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3238;
      end
      12'b110010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3239;
      end
      12'b110010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3240;
      end
      12'b110010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3241;
      end
      12'b110010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3242;
      end
      12'b110010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3243;
      end
      12'b110010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3244;
      end
      12'b110010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3245;
      end
      12'b110010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3246;
      end
      12'b110010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3247;
      end
      12'b110010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3248;
      end
      12'b110010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3249;
      end
      12'b110010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3250;
      end
      12'b110010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3251;
      end
      12'b110010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3252;
      end
      12'b110010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3253;
      end
      12'b110010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3254;
      end
      12'b110010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3255;
      end
      12'b110010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3256;
      end
      12'b110010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3257;
      end
      12'b110010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3258;
      end
      12'b110010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3259;
      end
      12'b110010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3260;
      end
      12'b110010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3261;
      end
      12'b110010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3262;
      end
      12'b110010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3263;
      end
      12'b110011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3264;
      end
      12'b110011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3265;
      end
      12'b110011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3266;
      end
      12'b110011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3267;
      end
      12'b110011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3268;
      end
      12'b110011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3269;
      end
      12'b110011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3270;
      end
      12'b110011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3271;
      end
      12'b110011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3272;
      end
      12'b110011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3273;
      end
      12'b110011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3274;
      end
      12'b110011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3275;
      end
      12'b110011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3276;
      end
      12'b110011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3277;
      end
      12'b110011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3278;
      end
      12'b110011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3279;
      end
      12'b110011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3280;
      end
      12'b110011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3281;
      end
      12'b110011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3282;
      end
      12'b110011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3283;
      end
      12'b110011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3284;
      end
      12'b110011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3285;
      end
      12'b110011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3286;
      end
      12'b110011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3287;
      end
      12'b110011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3288;
      end
      12'b110011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3289;
      end
      12'b110011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3290;
      end
      12'b110011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3291;
      end
      12'b110011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3292;
      end
      12'b110011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3293;
      end
      12'b110011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3294;
      end
      12'b110011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3295;
      end
      12'b110011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3296;
      end
      12'b110011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3297;
      end
      12'b110011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3298;
      end
      12'b110011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3299;
      end
      12'b110011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3300;
      end
      12'b110011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3301;
      end
      12'b110011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3302;
      end
      12'b110011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3303;
      end
      12'b110011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3304;
      end
      12'b110011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3305;
      end
      12'b110011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3306;
      end
      12'b110011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3307;
      end
      12'b110011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3308;
      end
      12'b110011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3309;
      end
      12'b110011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3310;
      end
      12'b110011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3311;
      end
      12'b110011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3312;
      end
      12'b110011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3313;
      end
      12'b110011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3314;
      end
      12'b110011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3315;
      end
      12'b110011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3316;
      end
      12'b110011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3317;
      end
      12'b110011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3318;
      end
      12'b110011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3319;
      end
      12'b110011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3320;
      end
      12'b110011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3321;
      end
      12'b110011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3322;
      end
      12'b110011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3323;
      end
      12'b110011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3324;
      end
      12'b110011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3325;
      end
      12'b110011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3326;
      end
      12'b110011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3327;
      end
      12'b110100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3328;
      end
      12'b110100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3329;
      end
      12'b110100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3330;
      end
      12'b110100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3331;
      end
      12'b110100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3332;
      end
      12'b110100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3333;
      end
      12'b110100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3334;
      end
      12'b110100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3335;
      end
      12'b110100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3336;
      end
      12'b110100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3337;
      end
      12'b110100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3338;
      end
      12'b110100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3339;
      end
      12'b110100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3340;
      end
      12'b110100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3341;
      end
      12'b110100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3342;
      end
      12'b110100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3343;
      end
      12'b110100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3344;
      end
      12'b110100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3345;
      end
      12'b110100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3346;
      end
      12'b110100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3347;
      end
      12'b110100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3348;
      end
      12'b110100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3349;
      end
      12'b110100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3350;
      end
      12'b110100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3351;
      end
      12'b110100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3352;
      end
      12'b110100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3353;
      end
      12'b110100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3354;
      end
      12'b110100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3355;
      end
      12'b110100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3356;
      end
      12'b110100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3357;
      end
      12'b110100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3358;
      end
      12'b110100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3359;
      end
      12'b110100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3360;
      end
      12'b110100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3361;
      end
      12'b110100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3362;
      end
      12'b110100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3363;
      end
      12'b110100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3364;
      end
      12'b110100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3365;
      end
      12'b110100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3366;
      end
      12'b110100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3367;
      end
      12'b110100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3368;
      end
      12'b110100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3369;
      end
      12'b110100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3370;
      end
      12'b110100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3371;
      end
      12'b110100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3372;
      end
      12'b110100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3373;
      end
      12'b110100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3374;
      end
      12'b110100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3375;
      end
      12'b110100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3376;
      end
      12'b110100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3377;
      end
      12'b110100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3378;
      end
      12'b110100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3379;
      end
      12'b110100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3380;
      end
      12'b110100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3381;
      end
      12'b110100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3382;
      end
      12'b110100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3383;
      end
      12'b110100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3384;
      end
      12'b110100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3385;
      end
      12'b110100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3386;
      end
      12'b110100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3387;
      end
      12'b110100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3388;
      end
      12'b110100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3389;
      end
      12'b110100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3390;
      end
      12'b110100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3391;
      end
      12'b110101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3392;
      end
      12'b110101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3393;
      end
      12'b110101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3394;
      end
      12'b110101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3395;
      end
      12'b110101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3396;
      end
      12'b110101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3397;
      end
      12'b110101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3398;
      end
      12'b110101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3399;
      end
      12'b110101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3400;
      end
      12'b110101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3401;
      end
      12'b110101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3402;
      end
      12'b110101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3403;
      end
      12'b110101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3404;
      end
      12'b110101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3405;
      end
      12'b110101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3406;
      end
      12'b110101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3407;
      end
      12'b110101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3408;
      end
      12'b110101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3409;
      end
      12'b110101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3410;
      end
      12'b110101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3411;
      end
      12'b110101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3412;
      end
      12'b110101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3413;
      end
      12'b110101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3414;
      end
      12'b110101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3415;
      end
      12'b110101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3416;
      end
      12'b110101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3417;
      end
      12'b110101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3418;
      end
      12'b110101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3419;
      end
      12'b110101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3420;
      end
      12'b110101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3421;
      end
      12'b110101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3422;
      end
      12'b110101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3423;
      end
      12'b110101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3424;
      end
      12'b110101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3425;
      end
      12'b110101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3426;
      end
      12'b110101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3427;
      end
      12'b110101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3428;
      end
      12'b110101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3429;
      end
      12'b110101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3430;
      end
      12'b110101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3431;
      end
      12'b110101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3432;
      end
      12'b110101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3433;
      end
      12'b110101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3434;
      end
      12'b110101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3435;
      end
      12'b110101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3436;
      end
      12'b110101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3437;
      end
      12'b110101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3438;
      end
      12'b110101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3439;
      end
      12'b110101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3440;
      end
      12'b110101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3441;
      end
      12'b110101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3442;
      end
      12'b110101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3443;
      end
      12'b110101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3444;
      end
      12'b110101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3445;
      end
      12'b110101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3446;
      end
      12'b110101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3447;
      end
      12'b110101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3448;
      end
      12'b110101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3449;
      end
      12'b110101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3450;
      end
      12'b110101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3451;
      end
      12'b110101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3452;
      end
      12'b110101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3453;
      end
      12'b110101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3454;
      end
      12'b110101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3455;
      end
      12'b110110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3456;
      end
      12'b110110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3457;
      end
      12'b110110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3458;
      end
      12'b110110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3459;
      end
      12'b110110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3460;
      end
      12'b110110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3461;
      end
      12'b110110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3462;
      end
      12'b110110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3463;
      end
      12'b110110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3464;
      end
      12'b110110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3465;
      end
      12'b110110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3466;
      end
      12'b110110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3467;
      end
      12'b110110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3468;
      end
      12'b110110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3469;
      end
      12'b110110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3470;
      end
      12'b110110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3471;
      end
      12'b110110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3472;
      end
      12'b110110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3473;
      end
      12'b110110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3474;
      end
      12'b110110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3475;
      end
      12'b110110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3476;
      end
      12'b110110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3477;
      end
      12'b110110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3478;
      end
      12'b110110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3479;
      end
      12'b110110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3480;
      end
      12'b110110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3481;
      end
      12'b110110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3482;
      end
      12'b110110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3483;
      end
      12'b110110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3484;
      end
      12'b110110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3485;
      end
      12'b110110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3486;
      end
      12'b110110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3487;
      end
      12'b110110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3488;
      end
      12'b110110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3489;
      end
      12'b110110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3490;
      end
      12'b110110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3491;
      end
      12'b110110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3492;
      end
      12'b110110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3493;
      end
      12'b110110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3494;
      end
      12'b110110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3495;
      end
      12'b110110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3496;
      end
      12'b110110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3497;
      end
      12'b110110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3498;
      end
      12'b110110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3499;
      end
      12'b110110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3500;
      end
      12'b110110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3501;
      end
      12'b110110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3502;
      end
      12'b110110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3503;
      end
      12'b110110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3504;
      end
      12'b110110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3505;
      end
      12'b110110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3506;
      end
      12'b110110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3507;
      end
      12'b110110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3508;
      end
      12'b110110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3509;
      end
      12'b110110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3510;
      end
      12'b110110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3511;
      end
      12'b110110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3512;
      end
      12'b110110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3513;
      end
      12'b110110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3514;
      end
      12'b110110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3515;
      end
      12'b110110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3516;
      end
      12'b110110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3517;
      end
      12'b110110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3518;
      end
      12'b110110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3519;
      end
      12'b110111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3520;
      end
      12'b110111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3521;
      end
      12'b110111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3522;
      end
      12'b110111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3523;
      end
      12'b110111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3524;
      end
      12'b110111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3525;
      end
      12'b110111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3526;
      end
      12'b110111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3527;
      end
      12'b110111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3528;
      end
      12'b110111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3529;
      end
      12'b110111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3530;
      end
      12'b110111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3531;
      end
      12'b110111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3532;
      end
      12'b110111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3533;
      end
      12'b110111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3534;
      end
      12'b110111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3535;
      end
      12'b110111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3536;
      end
      12'b110111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3537;
      end
      12'b110111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3538;
      end
      12'b110111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3539;
      end
      12'b110111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3540;
      end
      12'b110111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3541;
      end
      12'b110111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3542;
      end
      12'b110111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3543;
      end
      12'b110111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3544;
      end
      12'b110111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3545;
      end
      12'b110111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3546;
      end
      12'b110111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3547;
      end
      12'b110111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3548;
      end
      12'b110111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3549;
      end
      12'b110111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3550;
      end
      12'b110111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3551;
      end
      12'b110111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3552;
      end
      12'b110111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3553;
      end
      12'b110111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3554;
      end
      12'b110111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3555;
      end
      12'b110111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3556;
      end
      12'b110111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3557;
      end
      12'b110111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3558;
      end
      12'b110111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3559;
      end
      12'b110111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3560;
      end
      12'b110111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3561;
      end
      12'b110111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3562;
      end
      12'b110111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3563;
      end
      12'b110111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3564;
      end
      12'b110111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3565;
      end
      12'b110111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3566;
      end
      12'b110111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3567;
      end
      12'b110111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3568;
      end
      12'b110111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3569;
      end
      12'b110111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3570;
      end
      12'b110111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3571;
      end
      12'b110111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3572;
      end
      12'b110111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3573;
      end
      12'b110111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3574;
      end
      12'b110111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3575;
      end
      12'b110111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3576;
      end
      12'b110111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3577;
      end
      12'b110111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3578;
      end
      12'b110111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3579;
      end
      12'b110111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3580;
      end
      12'b110111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3581;
      end
      12'b110111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3582;
      end
      12'b110111111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3583;
      end
      12'b111000000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3584;
      end
      12'b111000000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3585;
      end
      12'b111000000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3586;
      end
      12'b111000000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3587;
      end
      12'b111000000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3588;
      end
      12'b111000000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3589;
      end
      12'b111000000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3590;
      end
      12'b111000000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3591;
      end
      12'b111000001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3592;
      end
      12'b111000001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3593;
      end
      12'b111000001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3594;
      end
      12'b111000001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3595;
      end
      12'b111000001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3596;
      end
      12'b111000001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3597;
      end
      12'b111000001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3598;
      end
      12'b111000001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3599;
      end
      12'b111000010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3600;
      end
      12'b111000010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3601;
      end
      12'b111000010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3602;
      end
      12'b111000010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3603;
      end
      12'b111000010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3604;
      end
      12'b111000010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3605;
      end
      12'b111000010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3606;
      end
      12'b111000010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3607;
      end
      12'b111000011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3608;
      end
      12'b111000011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3609;
      end
      12'b111000011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3610;
      end
      12'b111000011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3611;
      end
      12'b111000011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3612;
      end
      12'b111000011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3613;
      end
      12'b111000011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3614;
      end
      12'b111000011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3615;
      end
      12'b111000100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3616;
      end
      12'b111000100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3617;
      end
      12'b111000100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3618;
      end
      12'b111000100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3619;
      end
      12'b111000100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3620;
      end
      12'b111000100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3621;
      end
      12'b111000100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3622;
      end
      12'b111000100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3623;
      end
      12'b111000101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3624;
      end
      12'b111000101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3625;
      end
      12'b111000101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3626;
      end
      12'b111000101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3627;
      end
      12'b111000101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3628;
      end
      12'b111000101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3629;
      end
      12'b111000101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3630;
      end
      12'b111000101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3631;
      end
      12'b111000110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3632;
      end
      12'b111000110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3633;
      end
      12'b111000110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3634;
      end
      12'b111000110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3635;
      end
      12'b111000110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3636;
      end
      12'b111000110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3637;
      end
      12'b111000110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3638;
      end
      12'b111000110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3639;
      end
      12'b111000111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3640;
      end
      12'b111000111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3641;
      end
      12'b111000111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3642;
      end
      12'b111000111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3643;
      end
      12'b111000111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3644;
      end
      12'b111000111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3645;
      end
      12'b111000111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3646;
      end
      12'b111000111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3647;
      end
      12'b111001000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3648;
      end
      12'b111001000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3649;
      end
      12'b111001000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3650;
      end
      12'b111001000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3651;
      end
      12'b111001000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3652;
      end
      12'b111001000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3653;
      end
      12'b111001000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3654;
      end
      12'b111001000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3655;
      end
      12'b111001001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3656;
      end
      12'b111001001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3657;
      end
      12'b111001001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3658;
      end
      12'b111001001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3659;
      end
      12'b111001001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3660;
      end
      12'b111001001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3661;
      end
      12'b111001001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3662;
      end
      12'b111001001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3663;
      end
      12'b111001010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3664;
      end
      12'b111001010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3665;
      end
      12'b111001010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3666;
      end
      12'b111001010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3667;
      end
      12'b111001010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3668;
      end
      12'b111001010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3669;
      end
      12'b111001010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3670;
      end
      12'b111001010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3671;
      end
      12'b111001011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3672;
      end
      12'b111001011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3673;
      end
      12'b111001011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3674;
      end
      12'b111001011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3675;
      end
      12'b111001011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3676;
      end
      12'b111001011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3677;
      end
      12'b111001011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3678;
      end
      12'b111001011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3679;
      end
      12'b111001100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3680;
      end
      12'b111001100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3681;
      end
      12'b111001100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3682;
      end
      12'b111001100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3683;
      end
      12'b111001100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3684;
      end
      12'b111001100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3685;
      end
      12'b111001100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3686;
      end
      12'b111001100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3687;
      end
      12'b111001101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3688;
      end
      12'b111001101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3689;
      end
      12'b111001101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3690;
      end
      12'b111001101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3691;
      end
      12'b111001101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3692;
      end
      12'b111001101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3693;
      end
      12'b111001101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3694;
      end
      12'b111001101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3695;
      end
      12'b111001110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3696;
      end
      12'b111001110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3697;
      end
      12'b111001110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3698;
      end
      12'b111001110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3699;
      end
      12'b111001110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3700;
      end
      12'b111001110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3701;
      end
      12'b111001110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3702;
      end
      12'b111001110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3703;
      end
      12'b111001111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3704;
      end
      12'b111001111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3705;
      end
      12'b111001111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3706;
      end
      12'b111001111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3707;
      end
      12'b111001111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3708;
      end
      12'b111001111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3709;
      end
      12'b111001111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3710;
      end
      12'b111001111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3711;
      end
      12'b111010000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3712;
      end
      12'b111010000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3713;
      end
      12'b111010000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3714;
      end
      12'b111010000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3715;
      end
      12'b111010000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3716;
      end
      12'b111010000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3717;
      end
      12'b111010000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3718;
      end
      12'b111010000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3719;
      end
      12'b111010001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3720;
      end
      12'b111010001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3721;
      end
      12'b111010001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3722;
      end
      12'b111010001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3723;
      end
      12'b111010001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3724;
      end
      12'b111010001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3725;
      end
      12'b111010001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3726;
      end
      12'b111010001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3727;
      end
      12'b111010010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3728;
      end
      12'b111010010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3729;
      end
      12'b111010010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3730;
      end
      12'b111010010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3731;
      end
      12'b111010010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3732;
      end
      12'b111010010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3733;
      end
      12'b111010010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3734;
      end
      12'b111010010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3735;
      end
      12'b111010011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3736;
      end
      12'b111010011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3737;
      end
      12'b111010011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3738;
      end
      12'b111010011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3739;
      end
      12'b111010011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3740;
      end
      12'b111010011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3741;
      end
      12'b111010011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3742;
      end
      12'b111010011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3743;
      end
      12'b111010100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3744;
      end
      12'b111010100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3745;
      end
      12'b111010100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3746;
      end
      12'b111010100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3747;
      end
      12'b111010100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3748;
      end
      12'b111010100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3749;
      end
      12'b111010100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3750;
      end
      12'b111010100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3751;
      end
      12'b111010101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3752;
      end
      12'b111010101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3753;
      end
      12'b111010101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3754;
      end
      12'b111010101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3755;
      end
      12'b111010101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3756;
      end
      12'b111010101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3757;
      end
      12'b111010101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3758;
      end
      12'b111010101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3759;
      end
      12'b111010110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3760;
      end
      12'b111010110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3761;
      end
      12'b111010110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3762;
      end
      12'b111010110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3763;
      end
      12'b111010110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3764;
      end
      12'b111010110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3765;
      end
      12'b111010110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3766;
      end
      12'b111010110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3767;
      end
      12'b111010111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3768;
      end
      12'b111010111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3769;
      end
      12'b111010111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3770;
      end
      12'b111010111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3771;
      end
      12'b111010111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3772;
      end
      12'b111010111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3773;
      end
      12'b111010111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3774;
      end
      12'b111010111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3775;
      end
      12'b111011000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3776;
      end
      12'b111011000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3777;
      end
      12'b111011000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3778;
      end
      12'b111011000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3779;
      end
      12'b111011000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3780;
      end
      12'b111011000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3781;
      end
      12'b111011000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3782;
      end
      12'b111011000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3783;
      end
      12'b111011001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3784;
      end
      12'b111011001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3785;
      end
      12'b111011001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3786;
      end
      12'b111011001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3787;
      end
      12'b111011001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3788;
      end
      12'b111011001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3789;
      end
      12'b111011001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3790;
      end
      12'b111011001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3791;
      end
      12'b111011010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3792;
      end
      12'b111011010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3793;
      end
      12'b111011010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3794;
      end
      12'b111011010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3795;
      end
      12'b111011010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3796;
      end
      12'b111011010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3797;
      end
      12'b111011010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3798;
      end
      12'b111011010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3799;
      end
      12'b111011011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3800;
      end
      12'b111011011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3801;
      end
      12'b111011011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3802;
      end
      12'b111011011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3803;
      end
      12'b111011011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3804;
      end
      12'b111011011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3805;
      end
      12'b111011011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3806;
      end
      12'b111011011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3807;
      end
      12'b111011100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3808;
      end
      12'b111011100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3809;
      end
      12'b111011100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3810;
      end
      12'b111011100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3811;
      end
      12'b111011100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3812;
      end
      12'b111011100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3813;
      end
      12'b111011100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3814;
      end
      12'b111011100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3815;
      end
      12'b111011101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3816;
      end
      12'b111011101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3817;
      end
      12'b111011101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3818;
      end
      12'b111011101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3819;
      end
      12'b111011101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3820;
      end
      12'b111011101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3821;
      end
      12'b111011101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3822;
      end
      12'b111011101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3823;
      end
      12'b111011110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3824;
      end
      12'b111011110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3825;
      end
      12'b111011110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3826;
      end
      12'b111011110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3827;
      end
      12'b111011110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3828;
      end
      12'b111011110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3829;
      end
      12'b111011110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3830;
      end
      12'b111011110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3831;
      end
      12'b111011111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3832;
      end
      12'b111011111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3833;
      end
      12'b111011111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3834;
      end
      12'b111011111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3835;
      end
      12'b111011111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3836;
      end
      12'b111011111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3837;
      end
      12'b111011111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3838;
      end
      12'b111011111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3839;
      end
      12'b111100000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3840;
      end
      12'b111100000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3841;
      end
      12'b111100000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3842;
      end
      12'b111100000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3843;
      end
      12'b111100000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3844;
      end
      12'b111100000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3845;
      end
      12'b111100000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3846;
      end
      12'b111100000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3847;
      end
      12'b111100001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3848;
      end
      12'b111100001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3849;
      end
      12'b111100001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3850;
      end
      12'b111100001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3851;
      end
      12'b111100001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3852;
      end
      12'b111100001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3853;
      end
      12'b111100001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3854;
      end
      12'b111100001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3855;
      end
      12'b111100010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3856;
      end
      12'b111100010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3857;
      end
      12'b111100010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3858;
      end
      12'b111100010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3859;
      end
      12'b111100010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3860;
      end
      12'b111100010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3861;
      end
      12'b111100010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3862;
      end
      12'b111100010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3863;
      end
      12'b111100011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3864;
      end
      12'b111100011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3865;
      end
      12'b111100011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3866;
      end
      12'b111100011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3867;
      end
      12'b111100011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3868;
      end
      12'b111100011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3869;
      end
      12'b111100011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3870;
      end
      12'b111100011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3871;
      end
      12'b111100100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3872;
      end
      12'b111100100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3873;
      end
      12'b111100100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3874;
      end
      12'b111100100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3875;
      end
      12'b111100100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3876;
      end
      12'b111100100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3877;
      end
      12'b111100100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3878;
      end
      12'b111100100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3879;
      end
      12'b111100101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3880;
      end
      12'b111100101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3881;
      end
      12'b111100101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3882;
      end
      12'b111100101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3883;
      end
      12'b111100101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3884;
      end
      12'b111100101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3885;
      end
      12'b111100101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3886;
      end
      12'b111100101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3887;
      end
      12'b111100110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3888;
      end
      12'b111100110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3889;
      end
      12'b111100110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3890;
      end
      12'b111100110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3891;
      end
      12'b111100110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3892;
      end
      12'b111100110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3893;
      end
      12'b111100110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3894;
      end
      12'b111100110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3895;
      end
      12'b111100111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3896;
      end
      12'b111100111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3897;
      end
      12'b111100111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3898;
      end
      12'b111100111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3899;
      end
      12'b111100111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3900;
      end
      12'b111100111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3901;
      end
      12'b111100111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3902;
      end
      12'b111100111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3903;
      end
      12'b111101000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3904;
      end
      12'b111101000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3905;
      end
      12'b111101000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3906;
      end
      12'b111101000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3907;
      end
      12'b111101000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3908;
      end
      12'b111101000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3909;
      end
      12'b111101000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3910;
      end
      12'b111101000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3911;
      end
      12'b111101001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3912;
      end
      12'b111101001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3913;
      end
      12'b111101001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3914;
      end
      12'b111101001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3915;
      end
      12'b111101001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3916;
      end
      12'b111101001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3917;
      end
      12'b111101001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3918;
      end
      12'b111101001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3919;
      end
      12'b111101010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3920;
      end
      12'b111101010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3921;
      end
      12'b111101010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3922;
      end
      12'b111101010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3923;
      end
      12'b111101010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3924;
      end
      12'b111101010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3925;
      end
      12'b111101010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3926;
      end
      12'b111101010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3927;
      end
      12'b111101011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3928;
      end
      12'b111101011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3929;
      end
      12'b111101011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3930;
      end
      12'b111101011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3931;
      end
      12'b111101011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3932;
      end
      12'b111101011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3933;
      end
      12'b111101011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3934;
      end
      12'b111101011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3935;
      end
      12'b111101100000 : begin
        _zz_axiSignal_r_payload_data = regVec_3936;
      end
      12'b111101100001 : begin
        _zz_axiSignal_r_payload_data = regVec_3937;
      end
      12'b111101100010 : begin
        _zz_axiSignal_r_payload_data = regVec_3938;
      end
      12'b111101100011 : begin
        _zz_axiSignal_r_payload_data = regVec_3939;
      end
      12'b111101100100 : begin
        _zz_axiSignal_r_payload_data = regVec_3940;
      end
      12'b111101100101 : begin
        _zz_axiSignal_r_payload_data = regVec_3941;
      end
      12'b111101100110 : begin
        _zz_axiSignal_r_payload_data = regVec_3942;
      end
      12'b111101100111 : begin
        _zz_axiSignal_r_payload_data = regVec_3943;
      end
      12'b111101101000 : begin
        _zz_axiSignal_r_payload_data = regVec_3944;
      end
      12'b111101101001 : begin
        _zz_axiSignal_r_payload_data = regVec_3945;
      end
      12'b111101101010 : begin
        _zz_axiSignal_r_payload_data = regVec_3946;
      end
      12'b111101101011 : begin
        _zz_axiSignal_r_payload_data = regVec_3947;
      end
      12'b111101101100 : begin
        _zz_axiSignal_r_payload_data = regVec_3948;
      end
      12'b111101101101 : begin
        _zz_axiSignal_r_payload_data = regVec_3949;
      end
      12'b111101101110 : begin
        _zz_axiSignal_r_payload_data = regVec_3950;
      end
      12'b111101101111 : begin
        _zz_axiSignal_r_payload_data = regVec_3951;
      end
      12'b111101110000 : begin
        _zz_axiSignal_r_payload_data = regVec_3952;
      end
      12'b111101110001 : begin
        _zz_axiSignal_r_payload_data = regVec_3953;
      end
      12'b111101110010 : begin
        _zz_axiSignal_r_payload_data = regVec_3954;
      end
      12'b111101110011 : begin
        _zz_axiSignal_r_payload_data = regVec_3955;
      end
      12'b111101110100 : begin
        _zz_axiSignal_r_payload_data = regVec_3956;
      end
      12'b111101110101 : begin
        _zz_axiSignal_r_payload_data = regVec_3957;
      end
      12'b111101110110 : begin
        _zz_axiSignal_r_payload_data = regVec_3958;
      end
      12'b111101110111 : begin
        _zz_axiSignal_r_payload_data = regVec_3959;
      end
      12'b111101111000 : begin
        _zz_axiSignal_r_payload_data = regVec_3960;
      end
      12'b111101111001 : begin
        _zz_axiSignal_r_payload_data = regVec_3961;
      end
      12'b111101111010 : begin
        _zz_axiSignal_r_payload_data = regVec_3962;
      end
      12'b111101111011 : begin
        _zz_axiSignal_r_payload_data = regVec_3963;
      end
      12'b111101111100 : begin
        _zz_axiSignal_r_payload_data = regVec_3964;
      end
      12'b111101111101 : begin
        _zz_axiSignal_r_payload_data = regVec_3965;
      end
      12'b111101111110 : begin
        _zz_axiSignal_r_payload_data = regVec_3966;
      end
      12'b111101111111 : begin
        _zz_axiSignal_r_payload_data = regVec_3967;
      end
      12'b111110000000 : begin
        _zz_axiSignal_r_payload_data = regVec_3968;
      end
      12'b111110000001 : begin
        _zz_axiSignal_r_payload_data = regVec_3969;
      end
      12'b111110000010 : begin
        _zz_axiSignal_r_payload_data = regVec_3970;
      end
      12'b111110000011 : begin
        _zz_axiSignal_r_payload_data = regVec_3971;
      end
      12'b111110000100 : begin
        _zz_axiSignal_r_payload_data = regVec_3972;
      end
      12'b111110000101 : begin
        _zz_axiSignal_r_payload_data = regVec_3973;
      end
      12'b111110000110 : begin
        _zz_axiSignal_r_payload_data = regVec_3974;
      end
      12'b111110000111 : begin
        _zz_axiSignal_r_payload_data = regVec_3975;
      end
      12'b111110001000 : begin
        _zz_axiSignal_r_payload_data = regVec_3976;
      end
      12'b111110001001 : begin
        _zz_axiSignal_r_payload_data = regVec_3977;
      end
      12'b111110001010 : begin
        _zz_axiSignal_r_payload_data = regVec_3978;
      end
      12'b111110001011 : begin
        _zz_axiSignal_r_payload_data = regVec_3979;
      end
      12'b111110001100 : begin
        _zz_axiSignal_r_payload_data = regVec_3980;
      end
      12'b111110001101 : begin
        _zz_axiSignal_r_payload_data = regVec_3981;
      end
      12'b111110001110 : begin
        _zz_axiSignal_r_payload_data = regVec_3982;
      end
      12'b111110001111 : begin
        _zz_axiSignal_r_payload_data = regVec_3983;
      end
      12'b111110010000 : begin
        _zz_axiSignal_r_payload_data = regVec_3984;
      end
      12'b111110010001 : begin
        _zz_axiSignal_r_payload_data = regVec_3985;
      end
      12'b111110010010 : begin
        _zz_axiSignal_r_payload_data = regVec_3986;
      end
      12'b111110010011 : begin
        _zz_axiSignal_r_payload_data = regVec_3987;
      end
      12'b111110010100 : begin
        _zz_axiSignal_r_payload_data = regVec_3988;
      end
      12'b111110010101 : begin
        _zz_axiSignal_r_payload_data = regVec_3989;
      end
      12'b111110010110 : begin
        _zz_axiSignal_r_payload_data = regVec_3990;
      end
      12'b111110010111 : begin
        _zz_axiSignal_r_payload_data = regVec_3991;
      end
      12'b111110011000 : begin
        _zz_axiSignal_r_payload_data = regVec_3992;
      end
      12'b111110011001 : begin
        _zz_axiSignal_r_payload_data = regVec_3993;
      end
      12'b111110011010 : begin
        _zz_axiSignal_r_payload_data = regVec_3994;
      end
      12'b111110011011 : begin
        _zz_axiSignal_r_payload_data = regVec_3995;
      end
      12'b111110011100 : begin
        _zz_axiSignal_r_payload_data = regVec_3996;
      end
      12'b111110011101 : begin
        _zz_axiSignal_r_payload_data = regVec_3997;
      end
      12'b111110011110 : begin
        _zz_axiSignal_r_payload_data = regVec_3998;
      end
      12'b111110011111 : begin
        _zz_axiSignal_r_payload_data = regVec_3999;
      end
      12'b111110100000 : begin
        _zz_axiSignal_r_payload_data = regVec_4000;
      end
      12'b111110100001 : begin
        _zz_axiSignal_r_payload_data = regVec_4001;
      end
      12'b111110100010 : begin
        _zz_axiSignal_r_payload_data = regVec_4002;
      end
      12'b111110100011 : begin
        _zz_axiSignal_r_payload_data = regVec_4003;
      end
      12'b111110100100 : begin
        _zz_axiSignal_r_payload_data = regVec_4004;
      end
      12'b111110100101 : begin
        _zz_axiSignal_r_payload_data = regVec_4005;
      end
      12'b111110100110 : begin
        _zz_axiSignal_r_payload_data = regVec_4006;
      end
      12'b111110100111 : begin
        _zz_axiSignal_r_payload_data = regVec_4007;
      end
      12'b111110101000 : begin
        _zz_axiSignal_r_payload_data = regVec_4008;
      end
      12'b111110101001 : begin
        _zz_axiSignal_r_payload_data = regVec_4009;
      end
      12'b111110101010 : begin
        _zz_axiSignal_r_payload_data = regVec_4010;
      end
      12'b111110101011 : begin
        _zz_axiSignal_r_payload_data = regVec_4011;
      end
      12'b111110101100 : begin
        _zz_axiSignal_r_payload_data = regVec_4012;
      end
      12'b111110101101 : begin
        _zz_axiSignal_r_payload_data = regVec_4013;
      end
      12'b111110101110 : begin
        _zz_axiSignal_r_payload_data = regVec_4014;
      end
      12'b111110101111 : begin
        _zz_axiSignal_r_payload_data = regVec_4015;
      end
      12'b111110110000 : begin
        _zz_axiSignal_r_payload_data = regVec_4016;
      end
      12'b111110110001 : begin
        _zz_axiSignal_r_payload_data = regVec_4017;
      end
      12'b111110110010 : begin
        _zz_axiSignal_r_payload_data = regVec_4018;
      end
      12'b111110110011 : begin
        _zz_axiSignal_r_payload_data = regVec_4019;
      end
      12'b111110110100 : begin
        _zz_axiSignal_r_payload_data = regVec_4020;
      end
      12'b111110110101 : begin
        _zz_axiSignal_r_payload_data = regVec_4021;
      end
      12'b111110110110 : begin
        _zz_axiSignal_r_payload_data = regVec_4022;
      end
      12'b111110110111 : begin
        _zz_axiSignal_r_payload_data = regVec_4023;
      end
      12'b111110111000 : begin
        _zz_axiSignal_r_payload_data = regVec_4024;
      end
      12'b111110111001 : begin
        _zz_axiSignal_r_payload_data = regVec_4025;
      end
      12'b111110111010 : begin
        _zz_axiSignal_r_payload_data = regVec_4026;
      end
      12'b111110111011 : begin
        _zz_axiSignal_r_payload_data = regVec_4027;
      end
      12'b111110111100 : begin
        _zz_axiSignal_r_payload_data = regVec_4028;
      end
      12'b111110111101 : begin
        _zz_axiSignal_r_payload_data = regVec_4029;
      end
      12'b111110111110 : begin
        _zz_axiSignal_r_payload_data = regVec_4030;
      end
      12'b111110111111 : begin
        _zz_axiSignal_r_payload_data = regVec_4031;
      end
      12'b111111000000 : begin
        _zz_axiSignal_r_payload_data = regVec_4032;
      end
      12'b111111000001 : begin
        _zz_axiSignal_r_payload_data = regVec_4033;
      end
      12'b111111000010 : begin
        _zz_axiSignal_r_payload_data = regVec_4034;
      end
      12'b111111000011 : begin
        _zz_axiSignal_r_payload_data = regVec_4035;
      end
      12'b111111000100 : begin
        _zz_axiSignal_r_payload_data = regVec_4036;
      end
      12'b111111000101 : begin
        _zz_axiSignal_r_payload_data = regVec_4037;
      end
      12'b111111000110 : begin
        _zz_axiSignal_r_payload_data = regVec_4038;
      end
      12'b111111000111 : begin
        _zz_axiSignal_r_payload_data = regVec_4039;
      end
      12'b111111001000 : begin
        _zz_axiSignal_r_payload_data = regVec_4040;
      end
      12'b111111001001 : begin
        _zz_axiSignal_r_payload_data = regVec_4041;
      end
      12'b111111001010 : begin
        _zz_axiSignal_r_payload_data = regVec_4042;
      end
      12'b111111001011 : begin
        _zz_axiSignal_r_payload_data = regVec_4043;
      end
      12'b111111001100 : begin
        _zz_axiSignal_r_payload_data = regVec_4044;
      end
      12'b111111001101 : begin
        _zz_axiSignal_r_payload_data = regVec_4045;
      end
      12'b111111001110 : begin
        _zz_axiSignal_r_payload_data = regVec_4046;
      end
      12'b111111001111 : begin
        _zz_axiSignal_r_payload_data = regVec_4047;
      end
      12'b111111010000 : begin
        _zz_axiSignal_r_payload_data = regVec_4048;
      end
      12'b111111010001 : begin
        _zz_axiSignal_r_payload_data = regVec_4049;
      end
      12'b111111010010 : begin
        _zz_axiSignal_r_payload_data = regVec_4050;
      end
      12'b111111010011 : begin
        _zz_axiSignal_r_payload_data = regVec_4051;
      end
      12'b111111010100 : begin
        _zz_axiSignal_r_payload_data = regVec_4052;
      end
      12'b111111010101 : begin
        _zz_axiSignal_r_payload_data = regVec_4053;
      end
      12'b111111010110 : begin
        _zz_axiSignal_r_payload_data = regVec_4054;
      end
      12'b111111010111 : begin
        _zz_axiSignal_r_payload_data = regVec_4055;
      end
      12'b111111011000 : begin
        _zz_axiSignal_r_payload_data = regVec_4056;
      end
      12'b111111011001 : begin
        _zz_axiSignal_r_payload_data = regVec_4057;
      end
      12'b111111011010 : begin
        _zz_axiSignal_r_payload_data = regVec_4058;
      end
      12'b111111011011 : begin
        _zz_axiSignal_r_payload_data = regVec_4059;
      end
      12'b111111011100 : begin
        _zz_axiSignal_r_payload_data = regVec_4060;
      end
      12'b111111011101 : begin
        _zz_axiSignal_r_payload_data = regVec_4061;
      end
      12'b111111011110 : begin
        _zz_axiSignal_r_payload_data = regVec_4062;
      end
      12'b111111011111 : begin
        _zz_axiSignal_r_payload_data = regVec_4063;
      end
      12'b111111100000 : begin
        _zz_axiSignal_r_payload_data = regVec_4064;
      end
      12'b111111100001 : begin
        _zz_axiSignal_r_payload_data = regVec_4065;
      end
      12'b111111100010 : begin
        _zz_axiSignal_r_payload_data = regVec_4066;
      end
      12'b111111100011 : begin
        _zz_axiSignal_r_payload_data = regVec_4067;
      end
      12'b111111100100 : begin
        _zz_axiSignal_r_payload_data = regVec_4068;
      end
      12'b111111100101 : begin
        _zz_axiSignal_r_payload_data = regVec_4069;
      end
      12'b111111100110 : begin
        _zz_axiSignal_r_payload_data = regVec_4070;
      end
      12'b111111100111 : begin
        _zz_axiSignal_r_payload_data = regVec_4071;
      end
      12'b111111101000 : begin
        _zz_axiSignal_r_payload_data = regVec_4072;
      end
      12'b111111101001 : begin
        _zz_axiSignal_r_payload_data = regVec_4073;
      end
      12'b111111101010 : begin
        _zz_axiSignal_r_payload_data = regVec_4074;
      end
      12'b111111101011 : begin
        _zz_axiSignal_r_payload_data = regVec_4075;
      end
      12'b111111101100 : begin
        _zz_axiSignal_r_payload_data = regVec_4076;
      end
      12'b111111101101 : begin
        _zz_axiSignal_r_payload_data = regVec_4077;
      end
      12'b111111101110 : begin
        _zz_axiSignal_r_payload_data = regVec_4078;
      end
      12'b111111101111 : begin
        _zz_axiSignal_r_payload_data = regVec_4079;
      end
      12'b111111110000 : begin
        _zz_axiSignal_r_payload_data = regVec_4080;
      end
      12'b111111110001 : begin
        _zz_axiSignal_r_payload_data = regVec_4081;
      end
      12'b111111110010 : begin
        _zz_axiSignal_r_payload_data = regVec_4082;
      end
      12'b111111110011 : begin
        _zz_axiSignal_r_payload_data = regVec_4083;
      end
      12'b111111110100 : begin
        _zz_axiSignal_r_payload_data = regVec_4084;
      end
      12'b111111110101 : begin
        _zz_axiSignal_r_payload_data = regVec_4085;
      end
      12'b111111110110 : begin
        _zz_axiSignal_r_payload_data = regVec_4086;
      end
      12'b111111110111 : begin
        _zz_axiSignal_r_payload_data = regVec_4087;
      end
      12'b111111111000 : begin
        _zz_axiSignal_r_payload_data = regVec_4088;
      end
      12'b111111111001 : begin
        _zz_axiSignal_r_payload_data = regVec_4089;
      end
      12'b111111111010 : begin
        _zz_axiSignal_r_payload_data = regVec_4090;
      end
      12'b111111111011 : begin
        _zz_axiSignal_r_payload_data = regVec_4091;
      end
      12'b111111111100 : begin
        _zz_axiSignal_r_payload_data = regVec_4092;
      end
      12'b111111111101 : begin
        _zz_axiSignal_r_payload_data = regVec_4093;
      end
      12'b111111111110 : begin
        _zz_axiSignal_r_payload_data = regVec_4094;
      end
      default : begin
        _zz_axiSignal_r_payload_data = regVec_4095;
      end
    endcase
  end

  always @(*) begin
    case(Axi4Incr_wrapCase_1)
      2'b00 : begin
        _zz_Axi4Incr_result_1 = {Axi4Incr_base_1[11 : 1],Axi4Incr_baseIncr_1[0 : 0]};
      end
      2'b01 : begin
        _zz_Axi4Incr_result_1 = {Axi4Incr_base_1[11 : 2],Axi4Incr_baseIncr_1[1 : 0]};
      end
      2'b10 : begin
        _zz_Axi4Incr_result_1 = {Axi4Incr_base_1[11 : 3],Axi4Incr_baseIncr_1[2 : 0]};
      end
      default : begin
        _zz_Axi4Incr_result_1 = {Axi4Incr_base_1[11 : 4],Axi4Incr_baseIncr_1[3 : 0]};
      end
    endcase
  end

  always @(*) begin
    rFireCounter_willIncrement = 1'b0;
    if(when_Axi4_transmission_l174) begin
      rFireCounter_willIncrement = 1'b1;
    end
  end

  assign rFireCounter_willClear = 1'b0;
  assign rFireCounter_willOverflowIfInc = (rFireCounter_value == 13'h1000);
  assign rFireCounter_willOverflow = (rFireCounter_willOverflowIfInc && rFireCounter_willIncrement);
  always @(*) begin
    if(rFireCounter_willOverflow) begin
      rFireCounter_valueNext = 13'h0;
    end else begin
      rFireCounter_valueNext = (rFireCounter_value + _zz_rFireCounter_valueNext);
    end
    if(rFireCounter_willClear) begin
      rFireCounter_valueNext = 13'h0;
    end
  end

  assign bytePerWord = 1'b1;
  assign resetSignalValue = 1'b0;
  assign axiSignal_aw_ready = (updataAw && apstart);
  assign when_Axi4_transmission_l66 = (axiSignal_aw_valid && axiSignal_aw_ready);
  assign when_Axi4_transmission_l68 = (axiSignal_w_payload_last && (axiSignal_w_valid && axiSignal_w_ready));
  assign when_Axi4_transmission_l72 = (axiSignal_aw_valid && axiSignal_aw_ready);
  assign axiSignal_w_ready = (! updataAw);
  assign when_Axi4_transmission_l91 = (axiSignal_w_valid && axiSignal_w_ready);
  assign when_Axi4_transmission_l92 = 1'b1;
  assign _zz_1 = ({4095'd0,1'b1} <<< _zz__zz_1);
  assign _zz_regVec_0 = (axiSignal_w_payload_strb[0] ? axiSignal_w_payload_data[7 : 0] : _zz__zz_regVec_0);
  assign _zz_2 = ({4095'd0,1'b1} <<< regAwAddr);
  assign _zz_regVec_0_1 = (axiSignal_w_payload_strb[0] ? axiSignal_w_payload_data : _zz__zz_regVec_0_1_1);
  assign Axi4Incr_sizeValue = 1'b1;
  assign Axi4Incr_alignMask = 12'h0;
  assign Axi4Incr_base = (_zz_Axi4Incr_base & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(regAwLen)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (2'b00 + _zz_Axi4Incr_wrapCase);
  always @(*) begin
    case(regAwBrust)
      2'b00 : begin
        Axi4Incr_result = regAwAddr;
      end
      2'b10 : begin
        Axi4Incr_result = _zz_Axi4Incr_result;
      end
      default : begin
        Axi4Incr_result = Axi4Incr_baseIncr;
      end
    endcase
  end

  assign axiSignal_b_payload_id = 4'b0000;
  assign axiSignal_b_payload_resp = 2'b00;
  assign when_Axi4_transmission_l128 = (axiSignal_w_payload_last && (axiSignal_w_valid && axiSignal_w_ready));
  assign axiSignal_b_valid = writeSuccess;
  assign when_Axi4_transmission_l132 = (axiSignal_b_valid && axiSignal_b_ready);
  assign axiSignal_ar_ready = (updataAr && apstart);
  assign when_Axi4_transmission_l138 = (axiSignal_ar_valid && axiSignal_ar_ready);
  assign when_Axi4_transmission_l140 = (axiSignal_r_payload_last && (axiSignal_r_valid && axiSignal_r_ready));
  assign when_Axi4_transmission_l144 = (axiSignal_ar_valid && axiSignal_ar_ready);
  always @(*) begin
    if(axireset) begin
      axiSignal_r_valid = 1'b0;
    end else begin
      axiSignal_r_valid = ((! updataAr) && (! AwArConflict));
    end
  end

  assign axiSignal_r_payload_data[7 : 0] = _zz_axiSignal_r_payload_data;
  assign axiSignal_r_payload_id = 4'b0000;
  assign axiSignal_r_payload_resp = 2'b00;
  assign when_Axi4_transmission_l171 = (axiSignal_r_valid && axiSignal_r_ready);
  assign Axi4Incr_sizeValue_1 = 1'b1;
  assign Axi4Incr_alignMask_1 = 12'h0;
  assign Axi4Incr_base_1 = (_zz_Axi4Incr_base_1_1 & (~ Axi4Incr_alignMask_1));
  assign Axi4Incr_baseIncr_1 = (Axi4Incr_base_1 + _zz_Axi4Incr_baseIncr_1);
  always @(*) begin
    casez(regArLen)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase_1 = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase_1 = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase_1 = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase_1 = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase_1 = (2'b00 + _zz_Axi4Incr_wrapCase_1);
  always @(*) begin
    case(regArBrust)
      2'b00 : begin
        Axi4Incr_result_1 = regArAddr;
      end
      2'b10 : begin
        Axi4Incr_result_1 = _zz_Axi4Incr_result_1;
      end
      default : begin
        Axi4Incr_result_1 = Axi4Incr_baseIncr_1;
      end
    endcase
  end

  assign when_Axi4_transmission_l174 = (axiSignal_r_valid && axiSignal_r_ready);
  assign when_Axi4_transmission_l177 = ((rFireCounter_value == _zz_when_Axi4_transmission_l177) && (axiSignal_r_valid && axiSignal_r_ready));
  assign axiSignal_r_payload_last = (regLast && (axiSignal_r_valid && axiSignal_r_ready));
  assign when_Axi4_transmission_l182 = (((rFireCounter_value == _zz_when_Axi4_transmission_l182) && (regArLen != 8'h0)) && (axiSignal_r_valid && axiSignal_r_ready));
  assign when_Axi4_transmission_l184 = (regLast && axiSignal_r_payload_last);
  assign when_Axi4_transmission_l189 = (((axiSignal_aw_valid && axiSignal_aw_ready) && (axiSignal_ar_valid && axiSignal_ar_ready)) && (axiSignal_aw_payload_addr == axiSignal_ar_payload_addr));
  assign when_Axi4_transmission_l191 = ((AwArConflict && (axiSignal_b_valid && axiSignal_b_ready)) && (axiSignal_b_payload_resp == 2'b00));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      regVec_0 <= 8'h0;
      regVec_1 <= 8'h0;
      regVec_2 <= 8'h0;
      regVec_3 <= 8'h0;
      regVec_4 <= 8'h0;
      regVec_5 <= 8'h0;
      regVec_6 <= 8'h0;
      regVec_7 <= 8'h0;
      regVec_8 <= 8'h0;
      regVec_9 <= 8'h0;
      regVec_10 <= 8'h0;
      regVec_11 <= 8'h0;
      regVec_12 <= 8'h0;
      regVec_13 <= 8'h0;
      regVec_14 <= 8'h0;
      regVec_15 <= 8'h0;
      regVec_16 <= 8'h0;
      regVec_17 <= 8'h0;
      regVec_18 <= 8'h0;
      regVec_19 <= 8'h0;
      regVec_20 <= 8'h0;
      regVec_21 <= 8'h0;
      regVec_22 <= 8'h0;
      regVec_23 <= 8'h0;
      regVec_24 <= 8'h0;
      regVec_25 <= 8'h0;
      regVec_26 <= 8'h0;
      regVec_27 <= 8'h0;
      regVec_28 <= 8'h0;
      regVec_29 <= 8'h0;
      regVec_30 <= 8'h0;
      regVec_31 <= 8'h0;
      regVec_32 <= 8'h0;
      regVec_33 <= 8'h0;
      regVec_34 <= 8'h0;
      regVec_35 <= 8'h0;
      regVec_36 <= 8'h0;
      regVec_37 <= 8'h0;
      regVec_38 <= 8'h0;
      regVec_39 <= 8'h0;
      regVec_40 <= 8'h0;
      regVec_41 <= 8'h0;
      regVec_42 <= 8'h0;
      regVec_43 <= 8'h0;
      regVec_44 <= 8'h0;
      regVec_45 <= 8'h0;
      regVec_46 <= 8'h0;
      regVec_47 <= 8'h0;
      regVec_48 <= 8'h0;
      regVec_49 <= 8'h0;
      regVec_50 <= 8'h0;
      regVec_51 <= 8'h0;
      regVec_52 <= 8'h0;
      regVec_53 <= 8'h0;
      regVec_54 <= 8'h0;
      regVec_55 <= 8'h0;
      regVec_56 <= 8'h0;
      regVec_57 <= 8'h0;
      regVec_58 <= 8'h0;
      regVec_59 <= 8'h0;
      regVec_60 <= 8'h0;
      regVec_61 <= 8'h0;
      regVec_62 <= 8'h0;
      regVec_63 <= 8'h0;
      regVec_64 <= 8'h0;
      regVec_65 <= 8'h0;
      regVec_66 <= 8'h0;
      regVec_67 <= 8'h0;
      regVec_68 <= 8'h0;
      regVec_69 <= 8'h0;
      regVec_70 <= 8'h0;
      regVec_71 <= 8'h0;
      regVec_72 <= 8'h0;
      regVec_73 <= 8'h0;
      regVec_74 <= 8'h0;
      regVec_75 <= 8'h0;
      regVec_76 <= 8'h0;
      regVec_77 <= 8'h0;
      regVec_78 <= 8'h0;
      regVec_79 <= 8'h0;
      regVec_80 <= 8'h0;
      regVec_81 <= 8'h0;
      regVec_82 <= 8'h0;
      regVec_83 <= 8'h0;
      regVec_84 <= 8'h0;
      regVec_85 <= 8'h0;
      regVec_86 <= 8'h0;
      regVec_87 <= 8'h0;
      regVec_88 <= 8'h0;
      regVec_89 <= 8'h0;
      regVec_90 <= 8'h0;
      regVec_91 <= 8'h0;
      regVec_92 <= 8'h0;
      regVec_93 <= 8'h0;
      regVec_94 <= 8'h0;
      regVec_95 <= 8'h0;
      regVec_96 <= 8'h0;
      regVec_97 <= 8'h0;
      regVec_98 <= 8'h0;
      regVec_99 <= 8'h0;
      regVec_100 <= 8'h0;
      regVec_101 <= 8'h0;
      regVec_102 <= 8'h0;
      regVec_103 <= 8'h0;
      regVec_104 <= 8'h0;
      regVec_105 <= 8'h0;
      regVec_106 <= 8'h0;
      regVec_107 <= 8'h0;
      regVec_108 <= 8'h0;
      regVec_109 <= 8'h0;
      regVec_110 <= 8'h0;
      regVec_111 <= 8'h0;
      regVec_112 <= 8'h0;
      regVec_113 <= 8'h0;
      regVec_114 <= 8'h0;
      regVec_115 <= 8'h0;
      regVec_116 <= 8'h0;
      regVec_117 <= 8'h0;
      regVec_118 <= 8'h0;
      regVec_119 <= 8'h0;
      regVec_120 <= 8'h0;
      regVec_121 <= 8'h0;
      regVec_122 <= 8'h0;
      regVec_123 <= 8'h0;
      regVec_124 <= 8'h0;
      regVec_125 <= 8'h0;
      regVec_126 <= 8'h0;
      regVec_127 <= 8'h0;
      regVec_128 <= 8'h0;
      regVec_129 <= 8'h0;
      regVec_130 <= 8'h0;
      regVec_131 <= 8'h0;
      regVec_132 <= 8'h0;
      regVec_133 <= 8'h0;
      regVec_134 <= 8'h0;
      regVec_135 <= 8'h0;
      regVec_136 <= 8'h0;
      regVec_137 <= 8'h0;
      regVec_138 <= 8'h0;
      regVec_139 <= 8'h0;
      regVec_140 <= 8'h0;
      regVec_141 <= 8'h0;
      regVec_142 <= 8'h0;
      regVec_143 <= 8'h0;
      regVec_144 <= 8'h0;
      regVec_145 <= 8'h0;
      regVec_146 <= 8'h0;
      regVec_147 <= 8'h0;
      regVec_148 <= 8'h0;
      regVec_149 <= 8'h0;
      regVec_150 <= 8'h0;
      regVec_151 <= 8'h0;
      regVec_152 <= 8'h0;
      regVec_153 <= 8'h0;
      regVec_154 <= 8'h0;
      regVec_155 <= 8'h0;
      regVec_156 <= 8'h0;
      regVec_157 <= 8'h0;
      regVec_158 <= 8'h0;
      regVec_159 <= 8'h0;
      regVec_160 <= 8'h0;
      regVec_161 <= 8'h0;
      regVec_162 <= 8'h0;
      regVec_163 <= 8'h0;
      regVec_164 <= 8'h0;
      regVec_165 <= 8'h0;
      regVec_166 <= 8'h0;
      regVec_167 <= 8'h0;
      regVec_168 <= 8'h0;
      regVec_169 <= 8'h0;
      regVec_170 <= 8'h0;
      regVec_171 <= 8'h0;
      regVec_172 <= 8'h0;
      regVec_173 <= 8'h0;
      regVec_174 <= 8'h0;
      regVec_175 <= 8'h0;
      regVec_176 <= 8'h0;
      regVec_177 <= 8'h0;
      regVec_178 <= 8'h0;
      regVec_179 <= 8'h0;
      regVec_180 <= 8'h0;
      regVec_181 <= 8'h0;
      regVec_182 <= 8'h0;
      regVec_183 <= 8'h0;
      regVec_184 <= 8'h0;
      regVec_185 <= 8'h0;
      regVec_186 <= 8'h0;
      regVec_187 <= 8'h0;
      regVec_188 <= 8'h0;
      regVec_189 <= 8'h0;
      regVec_190 <= 8'h0;
      regVec_191 <= 8'h0;
      regVec_192 <= 8'h0;
      regVec_193 <= 8'h0;
      regVec_194 <= 8'h0;
      regVec_195 <= 8'h0;
      regVec_196 <= 8'h0;
      regVec_197 <= 8'h0;
      regVec_198 <= 8'h0;
      regVec_199 <= 8'h0;
      regVec_200 <= 8'h0;
      regVec_201 <= 8'h0;
      regVec_202 <= 8'h0;
      regVec_203 <= 8'h0;
      regVec_204 <= 8'h0;
      regVec_205 <= 8'h0;
      regVec_206 <= 8'h0;
      regVec_207 <= 8'h0;
      regVec_208 <= 8'h0;
      regVec_209 <= 8'h0;
      regVec_210 <= 8'h0;
      regVec_211 <= 8'h0;
      regVec_212 <= 8'h0;
      regVec_213 <= 8'h0;
      regVec_214 <= 8'h0;
      regVec_215 <= 8'h0;
      regVec_216 <= 8'h0;
      regVec_217 <= 8'h0;
      regVec_218 <= 8'h0;
      regVec_219 <= 8'h0;
      regVec_220 <= 8'h0;
      regVec_221 <= 8'h0;
      regVec_222 <= 8'h0;
      regVec_223 <= 8'h0;
      regVec_224 <= 8'h0;
      regVec_225 <= 8'h0;
      regVec_226 <= 8'h0;
      regVec_227 <= 8'h0;
      regVec_228 <= 8'h0;
      regVec_229 <= 8'h0;
      regVec_230 <= 8'h0;
      regVec_231 <= 8'h0;
      regVec_232 <= 8'h0;
      regVec_233 <= 8'h0;
      regVec_234 <= 8'h0;
      regVec_235 <= 8'h0;
      regVec_236 <= 8'h0;
      regVec_237 <= 8'h0;
      regVec_238 <= 8'h0;
      regVec_239 <= 8'h0;
      regVec_240 <= 8'h0;
      regVec_241 <= 8'h0;
      regVec_242 <= 8'h0;
      regVec_243 <= 8'h0;
      regVec_244 <= 8'h0;
      regVec_245 <= 8'h0;
      regVec_246 <= 8'h0;
      regVec_247 <= 8'h0;
      regVec_248 <= 8'h0;
      regVec_249 <= 8'h0;
      regVec_250 <= 8'h0;
      regVec_251 <= 8'h0;
      regVec_252 <= 8'h0;
      regVec_253 <= 8'h0;
      regVec_254 <= 8'h0;
      regVec_255 <= 8'h0;
      regVec_256 <= 8'h0;
      regVec_257 <= 8'h0;
      regVec_258 <= 8'h0;
      regVec_259 <= 8'h0;
      regVec_260 <= 8'h0;
      regVec_261 <= 8'h0;
      regVec_262 <= 8'h0;
      regVec_263 <= 8'h0;
      regVec_264 <= 8'h0;
      regVec_265 <= 8'h0;
      regVec_266 <= 8'h0;
      regVec_267 <= 8'h0;
      regVec_268 <= 8'h0;
      regVec_269 <= 8'h0;
      regVec_270 <= 8'h0;
      regVec_271 <= 8'h0;
      regVec_272 <= 8'h0;
      regVec_273 <= 8'h0;
      regVec_274 <= 8'h0;
      regVec_275 <= 8'h0;
      regVec_276 <= 8'h0;
      regVec_277 <= 8'h0;
      regVec_278 <= 8'h0;
      regVec_279 <= 8'h0;
      regVec_280 <= 8'h0;
      regVec_281 <= 8'h0;
      regVec_282 <= 8'h0;
      regVec_283 <= 8'h0;
      regVec_284 <= 8'h0;
      regVec_285 <= 8'h0;
      regVec_286 <= 8'h0;
      regVec_287 <= 8'h0;
      regVec_288 <= 8'h0;
      regVec_289 <= 8'h0;
      regVec_290 <= 8'h0;
      regVec_291 <= 8'h0;
      regVec_292 <= 8'h0;
      regVec_293 <= 8'h0;
      regVec_294 <= 8'h0;
      regVec_295 <= 8'h0;
      regVec_296 <= 8'h0;
      regVec_297 <= 8'h0;
      regVec_298 <= 8'h0;
      regVec_299 <= 8'h0;
      regVec_300 <= 8'h0;
      regVec_301 <= 8'h0;
      regVec_302 <= 8'h0;
      regVec_303 <= 8'h0;
      regVec_304 <= 8'h0;
      regVec_305 <= 8'h0;
      regVec_306 <= 8'h0;
      regVec_307 <= 8'h0;
      regVec_308 <= 8'h0;
      regVec_309 <= 8'h0;
      regVec_310 <= 8'h0;
      regVec_311 <= 8'h0;
      regVec_312 <= 8'h0;
      regVec_313 <= 8'h0;
      regVec_314 <= 8'h0;
      regVec_315 <= 8'h0;
      regVec_316 <= 8'h0;
      regVec_317 <= 8'h0;
      regVec_318 <= 8'h0;
      regVec_319 <= 8'h0;
      regVec_320 <= 8'h0;
      regVec_321 <= 8'h0;
      regVec_322 <= 8'h0;
      regVec_323 <= 8'h0;
      regVec_324 <= 8'h0;
      regVec_325 <= 8'h0;
      regVec_326 <= 8'h0;
      regVec_327 <= 8'h0;
      regVec_328 <= 8'h0;
      regVec_329 <= 8'h0;
      regVec_330 <= 8'h0;
      regVec_331 <= 8'h0;
      regVec_332 <= 8'h0;
      regVec_333 <= 8'h0;
      regVec_334 <= 8'h0;
      regVec_335 <= 8'h0;
      regVec_336 <= 8'h0;
      regVec_337 <= 8'h0;
      regVec_338 <= 8'h0;
      regVec_339 <= 8'h0;
      regVec_340 <= 8'h0;
      regVec_341 <= 8'h0;
      regVec_342 <= 8'h0;
      regVec_343 <= 8'h0;
      regVec_344 <= 8'h0;
      regVec_345 <= 8'h0;
      regVec_346 <= 8'h0;
      regVec_347 <= 8'h0;
      regVec_348 <= 8'h0;
      regVec_349 <= 8'h0;
      regVec_350 <= 8'h0;
      regVec_351 <= 8'h0;
      regVec_352 <= 8'h0;
      regVec_353 <= 8'h0;
      regVec_354 <= 8'h0;
      regVec_355 <= 8'h0;
      regVec_356 <= 8'h0;
      regVec_357 <= 8'h0;
      regVec_358 <= 8'h0;
      regVec_359 <= 8'h0;
      regVec_360 <= 8'h0;
      regVec_361 <= 8'h0;
      regVec_362 <= 8'h0;
      regVec_363 <= 8'h0;
      regVec_364 <= 8'h0;
      regVec_365 <= 8'h0;
      regVec_366 <= 8'h0;
      regVec_367 <= 8'h0;
      regVec_368 <= 8'h0;
      regVec_369 <= 8'h0;
      regVec_370 <= 8'h0;
      regVec_371 <= 8'h0;
      regVec_372 <= 8'h0;
      regVec_373 <= 8'h0;
      regVec_374 <= 8'h0;
      regVec_375 <= 8'h0;
      regVec_376 <= 8'h0;
      regVec_377 <= 8'h0;
      regVec_378 <= 8'h0;
      regVec_379 <= 8'h0;
      regVec_380 <= 8'h0;
      regVec_381 <= 8'h0;
      regVec_382 <= 8'h0;
      regVec_383 <= 8'h0;
      regVec_384 <= 8'h0;
      regVec_385 <= 8'h0;
      regVec_386 <= 8'h0;
      regVec_387 <= 8'h0;
      regVec_388 <= 8'h0;
      regVec_389 <= 8'h0;
      regVec_390 <= 8'h0;
      regVec_391 <= 8'h0;
      regVec_392 <= 8'h0;
      regVec_393 <= 8'h0;
      regVec_394 <= 8'h0;
      regVec_395 <= 8'h0;
      regVec_396 <= 8'h0;
      regVec_397 <= 8'h0;
      regVec_398 <= 8'h0;
      regVec_399 <= 8'h0;
      regVec_400 <= 8'h0;
      regVec_401 <= 8'h0;
      regVec_402 <= 8'h0;
      regVec_403 <= 8'h0;
      regVec_404 <= 8'h0;
      regVec_405 <= 8'h0;
      regVec_406 <= 8'h0;
      regVec_407 <= 8'h0;
      regVec_408 <= 8'h0;
      regVec_409 <= 8'h0;
      regVec_410 <= 8'h0;
      regVec_411 <= 8'h0;
      regVec_412 <= 8'h0;
      regVec_413 <= 8'h0;
      regVec_414 <= 8'h0;
      regVec_415 <= 8'h0;
      regVec_416 <= 8'h0;
      regVec_417 <= 8'h0;
      regVec_418 <= 8'h0;
      regVec_419 <= 8'h0;
      regVec_420 <= 8'h0;
      regVec_421 <= 8'h0;
      regVec_422 <= 8'h0;
      regVec_423 <= 8'h0;
      regVec_424 <= 8'h0;
      regVec_425 <= 8'h0;
      regVec_426 <= 8'h0;
      regVec_427 <= 8'h0;
      regVec_428 <= 8'h0;
      regVec_429 <= 8'h0;
      regVec_430 <= 8'h0;
      regVec_431 <= 8'h0;
      regVec_432 <= 8'h0;
      regVec_433 <= 8'h0;
      regVec_434 <= 8'h0;
      regVec_435 <= 8'h0;
      regVec_436 <= 8'h0;
      regVec_437 <= 8'h0;
      regVec_438 <= 8'h0;
      regVec_439 <= 8'h0;
      regVec_440 <= 8'h0;
      regVec_441 <= 8'h0;
      regVec_442 <= 8'h0;
      regVec_443 <= 8'h0;
      regVec_444 <= 8'h0;
      regVec_445 <= 8'h0;
      regVec_446 <= 8'h0;
      regVec_447 <= 8'h0;
      regVec_448 <= 8'h0;
      regVec_449 <= 8'h0;
      regVec_450 <= 8'h0;
      regVec_451 <= 8'h0;
      regVec_452 <= 8'h0;
      regVec_453 <= 8'h0;
      regVec_454 <= 8'h0;
      regVec_455 <= 8'h0;
      regVec_456 <= 8'h0;
      regVec_457 <= 8'h0;
      regVec_458 <= 8'h0;
      regVec_459 <= 8'h0;
      regVec_460 <= 8'h0;
      regVec_461 <= 8'h0;
      regVec_462 <= 8'h0;
      regVec_463 <= 8'h0;
      regVec_464 <= 8'h0;
      regVec_465 <= 8'h0;
      regVec_466 <= 8'h0;
      regVec_467 <= 8'h0;
      regVec_468 <= 8'h0;
      regVec_469 <= 8'h0;
      regVec_470 <= 8'h0;
      regVec_471 <= 8'h0;
      regVec_472 <= 8'h0;
      regVec_473 <= 8'h0;
      regVec_474 <= 8'h0;
      regVec_475 <= 8'h0;
      regVec_476 <= 8'h0;
      regVec_477 <= 8'h0;
      regVec_478 <= 8'h0;
      regVec_479 <= 8'h0;
      regVec_480 <= 8'h0;
      regVec_481 <= 8'h0;
      regVec_482 <= 8'h0;
      regVec_483 <= 8'h0;
      regVec_484 <= 8'h0;
      regVec_485 <= 8'h0;
      regVec_486 <= 8'h0;
      regVec_487 <= 8'h0;
      regVec_488 <= 8'h0;
      regVec_489 <= 8'h0;
      regVec_490 <= 8'h0;
      regVec_491 <= 8'h0;
      regVec_492 <= 8'h0;
      regVec_493 <= 8'h0;
      regVec_494 <= 8'h0;
      regVec_495 <= 8'h0;
      regVec_496 <= 8'h0;
      regVec_497 <= 8'h0;
      regVec_498 <= 8'h0;
      regVec_499 <= 8'h0;
      regVec_500 <= 8'h0;
      regVec_501 <= 8'h0;
      regVec_502 <= 8'h0;
      regVec_503 <= 8'h0;
      regVec_504 <= 8'h0;
      regVec_505 <= 8'h0;
      regVec_506 <= 8'h0;
      regVec_507 <= 8'h0;
      regVec_508 <= 8'h0;
      regVec_509 <= 8'h0;
      regVec_510 <= 8'h0;
      regVec_511 <= 8'h0;
      regVec_512 <= 8'h0;
      regVec_513 <= 8'h0;
      regVec_514 <= 8'h0;
      regVec_515 <= 8'h0;
      regVec_516 <= 8'h0;
      regVec_517 <= 8'h0;
      regVec_518 <= 8'h0;
      regVec_519 <= 8'h0;
      regVec_520 <= 8'h0;
      regVec_521 <= 8'h0;
      regVec_522 <= 8'h0;
      regVec_523 <= 8'h0;
      regVec_524 <= 8'h0;
      regVec_525 <= 8'h0;
      regVec_526 <= 8'h0;
      regVec_527 <= 8'h0;
      regVec_528 <= 8'h0;
      regVec_529 <= 8'h0;
      regVec_530 <= 8'h0;
      regVec_531 <= 8'h0;
      regVec_532 <= 8'h0;
      regVec_533 <= 8'h0;
      regVec_534 <= 8'h0;
      regVec_535 <= 8'h0;
      regVec_536 <= 8'h0;
      regVec_537 <= 8'h0;
      regVec_538 <= 8'h0;
      regVec_539 <= 8'h0;
      regVec_540 <= 8'h0;
      regVec_541 <= 8'h0;
      regVec_542 <= 8'h0;
      regVec_543 <= 8'h0;
      regVec_544 <= 8'h0;
      regVec_545 <= 8'h0;
      regVec_546 <= 8'h0;
      regVec_547 <= 8'h0;
      regVec_548 <= 8'h0;
      regVec_549 <= 8'h0;
      regVec_550 <= 8'h0;
      regVec_551 <= 8'h0;
      regVec_552 <= 8'h0;
      regVec_553 <= 8'h0;
      regVec_554 <= 8'h0;
      regVec_555 <= 8'h0;
      regVec_556 <= 8'h0;
      regVec_557 <= 8'h0;
      regVec_558 <= 8'h0;
      regVec_559 <= 8'h0;
      regVec_560 <= 8'h0;
      regVec_561 <= 8'h0;
      regVec_562 <= 8'h0;
      regVec_563 <= 8'h0;
      regVec_564 <= 8'h0;
      regVec_565 <= 8'h0;
      regVec_566 <= 8'h0;
      regVec_567 <= 8'h0;
      regVec_568 <= 8'h0;
      regVec_569 <= 8'h0;
      regVec_570 <= 8'h0;
      regVec_571 <= 8'h0;
      regVec_572 <= 8'h0;
      regVec_573 <= 8'h0;
      regVec_574 <= 8'h0;
      regVec_575 <= 8'h0;
      regVec_576 <= 8'h0;
      regVec_577 <= 8'h0;
      regVec_578 <= 8'h0;
      regVec_579 <= 8'h0;
      regVec_580 <= 8'h0;
      regVec_581 <= 8'h0;
      regVec_582 <= 8'h0;
      regVec_583 <= 8'h0;
      regVec_584 <= 8'h0;
      regVec_585 <= 8'h0;
      regVec_586 <= 8'h0;
      regVec_587 <= 8'h0;
      regVec_588 <= 8'h0;
      regVec_589 <= 8'h0;
      regVec_590 <= 8'h0;
      regVec_591 <= 8'h0;
      regVec_592 <= 8'h0;
      regVec_593 <= 8'h0;
      regVec_594 <= 8'h0;
      regVec_595 <= 8'h0;
      regVec_596 <= 8'h0;
      regVec_597 <= 8'h0;
      regVec_598 <= 8'h0;
      regVec_599 <= 8'h0;
      regVec_600 <= 8'h0;
      regVec_601 <= 8'h0;
      regVec_602 <= 8'h0;
      regVec_603 <= 8'h0;
      regVec_604 <= 8'h0;
      regVec_605 <= 8'h0;
      regVec_606 <= 8'h0;
      regVec_607 <= 8'h0;
      regVec_608 <= 8'h0;
      regVec_609 <= 8'h0;
      regVec_610 <= 8'h0;
      regVec_611 <= 8'h0;
      regVec_612 <= 8'h0;
      regVec_613 <= 8'h0;
      regVec_614 <= 8'h0;
      regVec_615 <= 8'h0;
      regVec_616 <= 8'h0;
      regVec_617 <= 8'h0;
      regVec_618 <= 8'h0;
      regVec_619 <= 8'h0;
      regVec_620 <= 8'h0;
      regVec_621 <= 8'h0;
      regVec_622 <= 8'h0;
      regVec_623 <= 8'h0;
      regVec_624 <= 8'h0;
      regVec_625 <= 8'h0;
      regVec_626 <= 8'h0;
      regVec_627 <= 8'h0;
      regVec_628 <= 8'h0;
      regVec_629 <= 8'h0;
      regVec_630 <= 8'h0;
      regVec_631 <= 8'h0;
      regVec_632 <= 8'h0;
      regVec_633 <= 8'h0;
      regVec_634 <= 8'h0;
      regVec_635 <= 8'h0;
      regVec_636 <= 8'h0;
      regVec_637 <= 8'h0;
      regVec_638 <= 8'h0;
      regVec_639 <= 8'h0;
      regVec_640 <= 8'h0;
      regVec_641 <= 8'h0;
      regVec_642 <= 8'h0;
      regVec_643 <= 8'h0;
      regVec_644 <= 8'h0;
      regVec_645 <= 8'h0;
      regVec_646 <= 8'h0;
      regVec_647 <= 8'h0;
      regVec_648 <= 8'h0;
      regVec_649 <= 8'h0;
      regVec_650 <= 8'h0;
      regVec_651 <= 8'h0;
      regVec_652 <= 8'h0;
      regVec_653 <= 8'h0;
      regVec_654 <= 8'h0;
      regVec_655 <= 8'h0;
      regVec_656 <= 8'h0;
      regVec_657 <= 8'h0;
      regVec_658 <= 8'h0;
      regVec_659 <= 8'h0;
      regVec_660 <= 8'h0;
      regVec_661 <= 8'h0;
      regVec_662 <= 8'h0;
      regVec_663 <= 8'h0;
      regVec_664 <= 8'h0;
      regVec_665 <= 8'h0;
      regVec_666 <= 8'h0;
      regVec_667 <= 8'h0;
      regVec_668 <= 8'h0;
      regVec_669 <= 8'h0;
      regVec_670 <= 8'h0;
      regVec_671 <= 8'h0;
      regVec_672 <= 8'h0;
      regVec_673 <= 8'h0;
      regVec_674 <= 8'h0;
      regVec_675 <= 8'h0;
      regVec_676 <= 8'h0;
      regVec_677 <= 8'h0;
      regVec_678 <= 8'h0;
      regVec_679 <= 8'h0;
      regVec_680 <= 8'h0;
      regVec_681 <= 8'h0;
      regVec_682 <= 8'h0;
      regVec_683 <= 8'h0;
      regVec_684 <= 8'h0;
      regVec_685 <= 8'h0;
      regVec_686 <= 8'h0;
      regVec_687 <= 8'h0;
      regVec_688 <= 8'h0;
      regVec_689 <= 8'h0;
      regVec_690 <= 8'h0;
      regVec_691 <= 8'h0;
      regVec_692 <= 8'h0;
      regVec_693 <= 8'h0;
      regVec_694 <= 8'h0;
      regVec_695 <= 8'h0;
      regVec_696 <= 8'h0;
      regVec_697 <= 8'h0;
      regVec_698 <= 8'h0;
      regVec_699 <= 8'h0;
      regVec_700 <= 8'h0;
      regVec_701 <= 8'h0;
      regVec_702 <= 8'h0;
      regVec_703 <= 8'h0;
      regVec_704 <= 8'h0;
      regVec_705 <= 8'h0;
      regVec_706 <= 8'h0;
      regVec_707 <= 8'h0;
      regVec_708 <= 8'h0;
      regVec_709 <= 8'h0;
      regVec_710 <= 8'h0;
      regVec_711 <= 8'h0;
      regVec_712 <= 8'h0;
      regVec_713 <= 8'h0;
      regVec_714 <= 8'h0;
      regVec_715 <= 8'h0;
      regVec_716 <= 8'h0;
      regVec_717 <= 8'h0;
      regVec_718 <= 8'h0;
      regVec_719 <= 8'h0;
      regVec_720 <= 8'h0;
      regVec_721 <= 8'h0;
      regVec_722 <= 8'h0;
      regVec_723 <= 8'h0;
      regVec_724 <= 8'h0;
      regVec_725 <= 8'h0;
      regVec_726 <= 8'h0;
      regVec_727 <= 8'h0;
      regVec_728 <= 8'h0;
      regVec_729 <= 8'h0;
      regVec_730 <= 8'h0;
      regVec_731 <= 8'h0;
      regVec_732 <= 8'h0;
      regVec_733 <= 8'h0;
      regVec_734 <= 8'h0;
      regVec_735 <= 8'h0;
      regVec_736 <= 8'h0;
      regVec_737 <= 8'h0;
      regVec_738 <= 8'h0;
      regVec_739 <= 8'h0;
      regVec_740 <= 8'h0;
      regVec_741 <= 8'h0;
      regVec_742 <= 8'h0;
      regVec_743 <= 8'h0;
      regVec_744 <= 8'h0;
      regVec_745 <= 8'h0;
      regVec_746 <= 8'h0;
      regVec_747 <= 8'h0;
      regVec_748 <= 8'h0;
      regVec_749 <= 8'h0;
      regVec_750 <= 8'h0;
      regVec_751 <= 8'h0;
      regVec_752 <= 8'h0;
      regVec_753 <= 8'h0;
      regVec_754 <= 8'h0;
      regVec_755 <= 8'h0;
      regVec_756 <= 8'h0;
      regVec_757 <= 8'h0;
      regVec_758 <= 8'h0;
      regVec_759 <= 8'h0;
      regVec_760 <= 8'h0;
      regVec_761 <= 8'h0;
      regVec_762 <= 8'h0;
      regVec_763 <= 8'h0;
      regVec_764 <= 8'h0;
      regVec_765 <= 8'h0;
      regVec_766 <= 8'h0;
      regVec_767 <= 8'h0;
      regVec_768 <= 8'h0;
      regVec_769 <= 8'h0;
      regVec_770 <= 8'h0;
      regVec_771 <= 8'h0;
      regVec_772 <= 8'h0;
      regVec_773 <= 8'h0;
      regVec_774 <= 8'h0;
      regVec_775 <= 8'h0;
      regVec_776 <= 8'h0;
      regVec_777 <= 8'h0;
      regVec_778 <= 8'h0;
      regVec_779 <= 8'h0;
      regVec_780 <= 8'h0;
      regVec_781 <= 8'h0;
      regVec_782 <= 8'h0;
      regVec_783 <= 8'h0;
      regVec_784 <= 8'h0;
      regVec_785 <= 8'h0;
      regVec_786 <= 8'h0;
      regVec_787 <= 8'h0;
      regVec_788 <= 8'h0;
      regVec_789 <= 8'h0;
      regVec_790 <= 8'h0;
      regVec_791 <= 8'h0;
      regVec_792 <= 8'h0;
      regVec_793 <= 8'h0;
      regVec_794 <= 8'h0;
      regVec_795 <= 8'h0;
      regVec_796 <= 8'h0;
      regVec_797 <= 8'h0;
      regVec_798 <= 8'h0;
      regVec_799 <= 8'h0;
      regVec_800 <= 8'h0;
      regVec_801 <= 8'h0;
      regVec_802 <= 8'h0;
      regVec_803 <= 8'h0;
      regVec_804 <= 8'h0;
      regVec_805 <= 8'h0;
      regVec_806 <= 8'h0;
      regVec_807 <= 8'h0;
      regVec_808 <= 8'h0;
      regVec_809 <= 8'h0;
      regVec_810 <= 8'h0;
      regVec_811 <= 8'h0;
      regVec_812 <= 8'h0;
      regVec_813 <= 8'h0;
      regVec_814 <= 8'h0;
      regVec_815 <= 8'h0;
      regVec_816 <= 8'h0;
      regVec_817 <= 8'h0;
      regVec_818 <= 8'h0;
      regVec_819 <= 8'h0;
      regVec_820 <= 8'h0;
      regVec_821 <= 8'h0;
      regVec_822 <= 8'h0;
      regVec_823 <= 8'h0;
      regVec_824 <= 8'h0;
      regVec_825 <= 8'h0;
      regVec_826 <= 8'h0;
      regVec_827 <= 8'h0;
      regVec_828 <= 8'h0;
      regVec_829 <= 8'h0;
      regVec_830 <= 8'h0;
      regVec_831 <= 8'h0;
      regVec_832 <= 8'h0;
      regVec_833 <= 8'h0;
      regVec_834 <= 8'h0;
      regVec_835 <= 8'h0;
      regVec_836 <= 8'h0;
      regVec_837 <= 8'h0;
      regVec_838 <= 8'h0;
      regVec_839 <= 8'h0;
      regVec_840 <= 8'h0;
      regVec_841 <= 8'h0;
      regVec_842 <= 8'h0;
      regVec_843 <= 8'h0;
      regVec_844 <= 8'h0;
      regVec_845 <= 8'h0;
      regVec_846 <= 8'h0;
      regVec_847 <= 8'h0;
      regVec_848 <= 8'h0;
      regVec_849 <= 8'h0;
      regVec_850 <= 8'h0;
      regVec_851 <= 8'h0;
      regVec_852 <= 8'h0;
      regVec_853 <= 8'h0;
      regVec_854 <= 8'h0;
      regVec_855 <= 8'h0;
      regVec_856 <= 8'h0;
      regVec_857 <= 8'h0;
      regVec_858 <= 8'h0;
      regVec_859 <= 8'h0;
      regVec_860 <= 8'h0;
      regVec_861 <= 8'h0;
      regVec_862 <= 8'h0;
      regVec_863 <= 8'h0;
      regVec_864 <= 8'h0;
      regVec_865 <= 8'h0;
      regVec_866 <= 8'h0;
      regVec_867 <= 8'h0;
      regVec_868 <= 8'h0;
      regVec_869 <= 8'h0;
      regVec_870 <= 8'h0;
      regVec_871 <= 8'h0;
      regVec_872 <= 8'h0;
      regVec_873 <= 8'h0;
      regVec_874 <= 8'h0;
      regVec_875 <= 8'h0;
      regVec_876 <= 8'h0;
      regVec_877 <= 8'h0;
      regVec_878 <= 8'h0;
      regVec_879 <= 8'h0;
      regVec_880 <= 8'h0;
      regVec_881 <= 8'h0;
      regVec_882 <= 8'h0;
      regVec_883 <= 8'h0;
      regVec_884 <= 8'h0;
      regVec_885 <= 8'h0;
      regVec_886 <= 8'h0;
      regVec_887 <= 8'h0;
      regVec_888 <= 8'h0;
      regVec_889 <= 8'h0;
      regVec_890 <= 8'h0;
      regVec_891 <= 8'h0;
      regVec_892 <= 8'h0;
      regVec_893 <= 8'h0;
      regVec_894 <= 8'h0;
      regVec_895 <= 8'h0;
      regVec_896 <= 8'h0;
      regVec_897 <= 8'h0;
      regVec_898 <= 8'h0;
      regVec_899 <= 8'h0;
      regVec_900 <= 8'h0;
      regVec_901 <= 8'h0;
      regVec_902 <= 8'h0;
      regVec_903 <= 8'h0;
      regVec_904 <= 8'h0;
      regVec_905 <= 8'h0;
      regVec_906 <= 8'h0;
      regVec_907 <= 8'h0;
      regVec_908 <= 8'h0;
      regVec_909 <= 8'h0;
      regVec_910 <= 8'h0;
      regVec_911 <= 8'h0;
      regVec_912 <= 8'h0;
      regVec_913 <= 8'h0;
      regVec_914 <= 8'h0;
      regVec_915 <= 8'h0;
      regVec_916 <= 8'h0;
      regVec_917 <= 8'h0;
      regVec_918 <= 8'h0;
      regVec_919 <= 8'h0;
      regVec_920 <= 8'h0;
      regVec_921 <= 8'h0;
      regVec_922 <= 8'h0;
      regVec_923 <= 8'h0;
      regVec_924 <= 8'h0;
      regVec_925 <= 8'h0;
      regVec_926 <= 8'h0;
      regVec_927 <= 8'h0;
      regVec_928 <= 8'h0;
      regVec_929 <= 8'h0;
      regVec_930 <= 8'h0;
      regVec_931 <= 8'h0;
      regVec_932 <= 8'h0;
      regVec_933 <= 8'h0;
      regVec_934 <= 8'h0;
      regVec_935 <= 8'h0;
      regVec_936 <= 8'h0;
      regVec_937 <= 8'h0;
      regVec_938 <= 8'h0;
      regVec_939 <= 8'h0;
      regVec_940 <= 8'h0;
      regVec_941 <= 8'h0;
      regVec_942 <= 8'h0;
      regVec_943 <= 8'h0;
      regVec_944 <= 8'h0;
      regVec_945 <= 8'h0;
      regVec_946 <= 8'h0;
      regVec_947 <= 8'h0;
      regVec_948 <= 8'h0;
      regVec_949 <= 8'h0;
      regVec_950 <= 8'h0;
      regVec_951 <= 8'h0;
      regVec_952 <= 8'h0;
      regVec_953 <= 8'h0;
      regVec_954 <= 8'h0;
      regVec_955 <= 8'h0;
      regVec_956 <= 8'h0;
      regVec_957 <= 8'h0;
      regVec_958 <= 8'h0;
      regVec_959 <= 8'h0;
      regVec_960 <= 8'h0;
      regVec_961 <= 8'h0;
      regVec_962 <= 8'h0;
      regVec_963 <= 8'h0;
      regVec_964 <= 8'h0;
      regVec_965 <= 8'h0;
      regVec_966 <= 8'h0;
      regVec_967 <= 8'h0;
      regVec_968 <= 8'h0;
      regVec_969 <= 8'h0;
      regVec_970 <= 8'h0;
      regVec_971 <= 8'h0;
      regVec_972 <= 8'h0;
      regVec_973 <= 8'h0;
      regVec_974 <= 8'h0;
      regVec_975 <= 8'h0;
      regVec_976 <= 8'h0;
      regVec_977 <= 8'h0;
      regVec_978 <= 8'h0;
      regVec_979 <= 8'h0;
      regVec_980 <= 8'h0;
      regVec_981 <= 8'h0;
      regVec_982 <= 8'h0;
      regVec_983 <= 8'h0;
      regVec_984 <= 8'h0;
      regVec_985 <= 8'h0;
      regVec_986 <= 8'h0;
      regVec_987 <= 8'h0;
      regVec_988 <= 8'h0;
      regVec_989 <= 8'h0;
      regVec_990 <= 8'h0;
      regVec_991 <= 8'h0;
      regVec_992 <= 8'h0;
      regVec_993 <= 8'h0;
      regVec_994 <= 8'h0;
      regVec_995 <= 8'h0;
      regVec_996 <= 8'h0;
      regVec_997 <= 8'h0;
      regVec_998 <= 8'h0;
      regVec_999 <= 8'h0;
      regVec_1000 <= 8'h0;
      regVec_1001 <= 8'h0;
      regVec_1002 <= 8'h0;
      regVec_1003 <= 8'h0;
      regVec_1004 <= 8'h0;
      regVec_1005 <= 8'h0;
      regVec_1006 <= 8'h0;
      regVec_1007 <= 8'h0;
      regVec_1008 <= 8'h0;
      regVec_1009 <= 8'h0;
      regVec_1010 <= 8'h0;
      regVec_1011 <= 8'h0;
      regVec_1012 <= 8'h0;
      regVec_1013 <= 8'h0;
      regVec_1014 <= 8'h0;
      regVec_1015 <= 8'h0;
      regVec_1016 <= 8'h0;
      regVec_1017 <= 8'h0;
      regVec_1018 <= 8'h0;
      regVec_1019 <= 8'h0;
      regVec_1020 <= 8'h0;
      regVec_1021 <= 8'h0;
      regVec_1022 <= 8'h0;
      regVec_1023 <= 8'h0;
      regVec_1024 <= 8'h0;
      regVec_1025 <= 8'h0;
      regVec_1026 <= 8'h0;
      regVec_1027 <= 8'h0;
      regVec_1028 <= 8'h0;
      regVec_1029 <= 8'h0;
      regVec_1030 <= 8'h0;
      regVec_1031 <= 8'h0;
      regVec_1032 <= 8'h0;
      regVec_1033 <= 8'h0;
      regVec_1034 <= 8'h0;
      regVec_1035 <= 8'h0;
      regVec_1036 <= 8'h0;
      regVec_1037 <= 8'h0;
      regVec_1038 <= 8'h0;
      regVec_1039 <= 8'h0;
      regVec_1040 <= 8'h0;
      regVec_1041 <= 8'h0;
      regVec_1042 <= 8'h0;
      regVec_1043 <= 8'h0;
      regVec_1044 <= 8'h0;
      regVec_1045 <= 8'h0;
      regVec_1046 <= 8'h0;
      regVec_1047 <= 8'h0;
      regVec_1048 <= 8'h0;
      regVec_1049 <= 8'h0;
      regVec_1050 <= 8'h0;
      regVec_1051 <= 8'h0;
      regVec_1052 <= 8'h0;
      regVec_1053 <= 8'h0;
      regVec_1054 <= 8'h0;
      regVec_1055 <= 8'h0;
      regVec_1056 <= 8'h0;
      regVec_1057 <= 8'h0;
      regVec_1058 <= 8'h0;
      regVec_1059 <= 8'h0;
      regVec_1060 <= 8'h0;
      regVec_1061 <= 8'h0;
      regVec_1062 <= 8'h0;
      regVec_1063 <= 8'h0;
      regVec_1064 <= 8'h0;
      regVec_1065 <= 8'h0;
      regVec_1066 <= 8'h0;
      regVec_1067 <= 8'h0;
      regVec_1068 <= 8'h0;
      regVec_1069 <= 8'h0;
      regVec_1070 <= 8'h0;
      regVec_1071 <= 8'h0;
      regVec_1072 <= 8'h0;
      regVec_1073 <= 8'h0;
      regVec_1074 <= 8'h0;
      regVec_1075 <= 8'h0;
      regVec_1076 <= 8'h0;
      regVec_1077 <= 8'h0;
      regVec_1078 <= 8'h0;
      regVec_1079 <= 8'h0;
      regVec_1080 <= 8'h0;
      regVec_1081 <= 8'h0;
      regVec_1082 <= 8'h0;
      regVec_1083 <= 8'h0;
      regVec_1084 <= 8'h0;
      regVec_1085 <= 8'h0;
      regVec_1086 <= 8'h0;
      regVec_1087 <= 8'h0;
      regVec_1088 <= 8'h0;
      regVec_1089 <= 8'h0;
      regVec_1090 <= 8'h0;
      regVec_1091 <= 8'h0;
      regVec_1092 <= 8'h0;
      regVec_1093 <= 8'h0;
      regVec_1094 <= 8'h0;
      regVec_1095 <= 8'h0;
      regVec_1096 <= 8'h0;
      regVec_1097 <= 8'h0;
      regVec_1098 <= 8'h0;
      regVec_1099 <= 8'h0;
      regVec_1100 <= 8'h0;
      regVec_1101 <= 8'h0;
      regVec_1102 <= 8'h0;
      regVec_1103 <= 8'h0;
      regVec_1104 <= 8'h0;
      regVec_1105 <= 8'h0;
      regVec_1106 <= 8'h0;
      regVec_1107 <= 8'h0;
      regVec_1108 <= 8'h0;
      regVec_1109 <= 8'h0;
      regVec_1110 <= 8'h0;
      regVec_1111 <= 8'h0;
      regVec_1112 <= 8'h0;
      regVec_1113 <= 8'h0;
      regVec_1114 <= 8'h0;
      regVec_1115 <= 8'h0;
      regVec_1116 <= 8'h0;
      regVec_1117 <= 8'h0;
      regVec_1118 <= 8'h0;
      regVec_1119 <= 8'h0;
      regVec_1120 <= 8'h0;
      regVec_1121 <= 8'h0;
      regVec_1122 <= 8'h0;
      regVec_1123 <= 8'h0;
      regVec_1124 <= 8'h0;
      regVec_1125 <= 8'h0;
      regVec_1126 <= 8'h0;
      regVec_1127 <= 8'h0;
      regVec_1128 <= 8'h0;
      regVec_1129 <= 8'h0;
      regVec_1130 <= 8'h0;
      regVec_1131 <= 8'h0;
      regVec_1132 <= 8'h0;
      regVec_1133 <= 8'h0;
      regVec_1134 <= 8'h0;
      regVec_1135 <= 8'h0;
      regVec_1136 <= 8'h0;
      regVec_1137 <= 8'h0;
      regVec_1138 <= 8'h0;
      regVec_1139 <= 8'h0;
      regVec_1140 <= 8'h0;
      regVec_1141 <= 8'h0;
      regVec_1142 <= 8'h0;
      regVec_1143 <= 8'h0;
      regVec_1144 <= 8'h0;
      regVec_1145 <= 8'h0;
      regVec_1146 <= 8'h0;
      regVec_1147 <= 8'h0;
      regVec_1148 <= 8'h0;
      regVec_1149 <= 8'h0;
      regVec_1150 <= 8'h0;
      regVec_1151 <= 8'h0;
      regVec_1152 <= 8'h0;
      regVec_1153 <= 8'h0;
      regVec_1154 <= 8'h0;
      regVec_1155 <= 8'h0;
      regVec_1156 <= 8'h0;
      regVec_1157 <= 8'h0;
      regVec_1158 <= 8'h0;
      regVec_1159 <= 8'h0;
      regVec_1160 <= 8'h0;
      regVec_1161 <= 8'h0;
      regVec_1162 <= 8'h0;
      regVec_1163 <= 8'h0;
      regVec_1164 <= 8'h0;
      regVec_1165 <= 8'h0;
      regVec_1166 <= 8'h0;
      regVec_1167 <= 8'h0;
      regVec_1168 <= 8'h0;
      regVec_1169 <= 8'h0;
      regVec_1170 <= 8'h0;
      regVec_1171 <= 8'h0;
      regVec_1172 <= 8'h0;
      regVec_1173 <= 8'h0;
      regVec_1174 <= 8'h0;
      regVec_1175 <= 8'h0;
      regVec_1176 <= 8'h0;
      regVec_1177 <= 8'h0;
      regVec_1178 <= 8'h0;
      regVec_1179 <= 8'h0;
      regVec_1180 <= 8'h0;
      regVec_1181 <= 8'h0;
      regVec_1182 <= 8'h0;
      regVec_1183 <= 8'h0;
      regVec_1184 <= 8'h0;
      regVec_1185 <= 8'h0;
      regVec_1186 <= 8'h0;
      regVec_1187 <= 8'h0;
      regVec_1188 <= 8'h0;
      regVec_1189 <= 8'h0;
      regVec_1190 <= 8'h0;
      regVec_1191 <= 8'h0;
      regVec_1192 <= 8'h0;
      regVec_1193 <= 8'h0;
      regVec_1194 <= 8'h0;
      regVec_1195 <= 8'h0;
      regVec_1196 <= 8'h0;
      regVec_1197 <= 8'h0;
      regVec_1198 <= 8'h0;
      regVec_1199 <= 8'h0;
      regVec_1200 <= 8'h0;
      regVec_1201 <= 8'h0;
      regVec_1202 <= 8'h0;
      regVec_1203 <= 8'h0;
      regVec_1204 <= 8'h0;
      regVec_1205 <= 8'h0;
      regVec_1206 <= 8'h0;
      regVec_1207 <= 8'h0;
      regVec_1208 <= 8'h0;
      regVec_1209 <= 8'h0;
      regVec_1210 <= 8'h0;
      regVec_1211 <= 8'h0;
      regVec_1212 <= 8'h0;
      regVec_1213 <= 8'h0;
      regVec_1214 <= 8'h0;
      regVec_1215 <= 8'h0;
      regVec_1216 <= 8'h0;
      regVec_1217 <= 8'h0;
      regVec_1218 <= 8'h0;
      regVec_1219 <= 8'h0;
      regVec_1220 <= 8'h0;
      regVec_1221 <= 8'h0;
      regVec_1222 <= 8'h0;
      regVec_1223 <= 8'h0;
      regVec_1224 <= 8'h0;
      regVec_1225 <= 8'h0;
      regVec_1226 <= 8'h0;
      regVec_1227 <= 8'h0;
      regVec_1228 <= 8'h0;
      regVec_1229 <= 8'h0;
      regVec_1230 <= 8'h0;
      regVec_1231 <= 8'h0;
      regVec_1232 <= 8'h0;
      regVec_1233 <= 8'h0;
      regVec_1234 <= 8'h0;
      regVec_1235 <= 8'h0;
      regVec_1236 <= 8'h0;
      regVec_1237 <= 8'h0;
      regVec_1238 <= 8'h0;
      regVec_1239 <= 8'h0;
      regVec_1240 <= 8'h0;
      regVec_1241 <= 8'h0;
      regVec_1242 <= 8'h0;
      regVec_1243 <= 8'h0;
      regVec_1244 <= 8'h0;
      regVec_1245 <= 8'h0;
      regVec_1246 <= 8'h0;
      regVec_1247 <= 8'h0;
      regVec_1248 <= 8'h0;
      regVec_1249 <= 8'h0;
      regVec_1250 <= 8'h0;
      regVec_1251 <= 8'h0;
      regVec_1252 <= 8'h0;
      regVec_1253 <= 8'h0;
      regVec_1254 <= 8'h0;
      regVec_1255 <= 8'h0;
      regVec_1256 <= 8'h0;
      regVec_1257 <= 8'h0;
      regVec_1258 <= 8'h0;
      regVec_1259 <= 8'h0;
      regVec_1260 <= 8'h0;
      regVec_1261 <= 8'h0;
      regVec_1262 <= 8'h0;
      regVec_1263 <= 8'h0;
      regVec_1264 <= 8'h0;
      regVec_1265 <= 8'h0;
      regVec_1266 <= 8'h0;
      regVec_1267 <= 8'h0;
      regVec_1268 <= 8'h0;
      regVec_1269 <= 8'h0;
      regVec_1270 <= 8'h0;
      regVec_1271 <= 8'h0;
      regVec_1272 <= 8'h0;
      regVec_1273 <= 8'h0;
      regVec_1274 <= 8'h0;
      regVec_1275 <= 8'h0;
      regVec_1276 <= 8'h0;
      regVec_1277 <= 8'h0;
      regVec_1278 <= 8'h0;
      regVec_1279 <= 8'h0;
      regVec_1280 <= 8'h0;
      regVec_1281 <= 8'h0;
      regVec_1282 <= 8'h0;
      regVec_1283 <= 8'h0;
      regVec_1284 <= 8'h0;
      regVec_1285 <= 8'h0;
      regVec_1286 <= 8'h0;
      regVec_1287 <= 8'h0;
      regVec_1288 <= 8'h0;
      regVec_1289 <= 8'h0;
      regVec_1290 <= 8'h0;
      regVec_1291 <= 8'h0;
      regVec_1292 <= 8'h0;
      regVec_1293 <= 8'h0;
      regVec_1294 <= 8'h0;
      regVec_1295 <= 8'h0;
      regVec_1296 <= 8'h0;
      regVec_1297 <= 8'h0;
      regVec_1298 <= 8'h0;
      regVec_1299 <= 8'h0;
      regVec_1300 <= 8'h0;
      regVec_1301 <= 8'h0;
      regVec_1302 <= 8'h0;
      regVec_1303 <= 8'h0;
      regVec_1304 <= 8'h0;
      regVec_1305 <= 8'h0;
      regVec_1306 <= 8'h0;
      regVec_1307 <= 8'h0;
      regVec_1308 <= 8'h0;
      regVec_1309 <= 8'h0;
      regVec_1310 <= 8'h0;
      regVec_1311 <= 8'h0;
      regVec_1312 <= 8'h0;
      regVec_1313 <= 8'h0;
      regVec_1314 <= 8'h0;
      regVec_1315 <= 8'h0;
      regVec_1316 <= 8'h0;
      regVec_1317 <= 8'h0;
      regVec_1318 <= 8'h0;
      regVec_1319 <= 8'h0;
      regVec_1320 <= 8'h0;
      regVec_1321 <= 8'h0;
      regVec_1322 <= 8'h0;
      regVec_1323 <= 8'h0;
      regVec_1324 <= 8'h0;
      regVec_1325 <= 8'h0;
      regVec_1326 <= 8'h0;
      regVec_1327 <= 8'h0;
      regVec_1328 <= 8'h0;
      regVec_1329 <= 8'h0;
      regVec_1330 <= 8'h0;
      regVec_1331 <= 8'h0;
      regVec_1332 <= 8'h0;
      regVec_1333 <= 8'h0;
      regVec_1334 <= 8'h0;
      regVec_1335 <= 8'h0;
      regVec_1336 <= 8'h0;
      regVec_1337 <= 8'h0;
      regVec_1338 <= 8'h0;
      regVec_1339 <= 8'h0;
      regVec_1340 <= 8'h0;
      regVec_1341 <= 8'h0;
      regVec_1342 <= 8'h0;
      regVec_1343 <= 8'h0;
      regVec_1344 <= 8'h0;
      regVec_1345 <= 8'h0;
      regVec_1346 <= 8'h0;
      regVec_1347 <= 8'h0;
      regVec_1348 <= 8'h0;
      regVec_1349 <= 8'h0;
      regVec_1350 <= 8'h0;
      regVec_1351 <= 8'h0;
      regVec_1352 <= 8'h0;
      regVec_1353 <= 8'h0;
      regVec_1354 <= 8'h0;
      regVec_1355 <= 8'h0;
      regVec_1356 <= 8'h0;
      regVec_1357 <= 8'h0;
      regVec_1358 <= 8'h0;
      regVec_1359 <= 8'h0;
      regVec_1360 <= 8'h0;
      regVec_1361 <= 8'h0;
      regVec_1362 <= 8'h0;
      regVec_1363 <= 8'h0;
      regVec_1364 <= 8'h0;
      regVec_1365 <= 8'h0;
      regVec_1366 <= 8'h0;
      regVec_1367 <= 8'h0;
      regVec_1368 <= 8'h0;
      regVec_1369 <= 8'h0;
      regVec_1370 <= 8'h0;
      regVec_1371 <= 8'h0;
      regVec_1372 <= 8'h0;
      regVec_1373 <= 8'h0;
      regVec_1374 <= 8'h0;
      regVec_1375 <= 8'h0;
      regVec_1376 <= 8'h0;
      regVec_1377 <= 8'h0;
      regVec_1378 <= 8'h0;
      regVec_1379 <= 8'h0;
      regVec_1380 <= 8'h0;
      regVec_1381 <= 8'h0;
      regVec_1382 <= 8'h0;
      regVec_1383 <= 8'h0;
      regVec_1384 <= 8'h0;
      regVec_1385 <= 8'h0;
      regVec_1386 <= 8'h0;
      regVec_1387 <= 8'h0;
      regVec_1388 <= 8'h0;
      regVec_1389 <= 8'h0;
      regVec_1390 <= 8'h0;
      regVec_1391 <= 8'h0;
      regVec_1392 <= 8'h0;
      regVec_1393 <= 8'h0;
      regVec_1394 <= 8'h0;
      regVec_1395 <= 8'h0;
      regVec_1396 <= 8'h0;
      regVec_1397 <= 8'h0;
      regVec_1398 <= 8'h0;
      regVec_1399 <= 8'h0;
      regVec_1400 <= 8'h0;
      regVec_1401 <= 8'h0;
      regVec_1402 <= 8'h0;
      regVec_1403 <= 8'h0;
      regVec_1404 <= 8'h0;
      regVec_1405 <= 8'h0;
      regVec_1406 <= 8'h0;
      regVec_1407 <= 8'h0;
      regVec_1408 <= 8'h0;
      regVec_1409 <= 8'h0;
      regVec_1410 <= 8'h0;
      regVec_1411 <= 8'h0;
      regVec_1412 <= 8'h0;
      regVec_1413 <= 8'h0;
      regVec_1414 <= 8'h0;
      regVec_1415 <= 8'h0;
      regVec_1416 <= 8'h0;
      regVec_1417 <= 8'h0;
      regVec_1418 <= 8'h0;
      regVec_1419 <= 8'h0;
      regVec_1420 <= 8'h0;
      regVec_1421 <= 8'h0;
      regVec_1422 <= 8'h0;
      regVec_1423 <= 8'h0;
      regVec_1424 <= 8'h0;
      regVec_1425 <= 8'h0;
      regVec_1426 <= 8'h0;
      regVec_1427 <= 8'h0;
      regVec_1428 <= 8'h0;
      regVec_1429 <= 8'h0;
      regVec_1430 <= 8'h0;
      regVec_1431 <= 8'h0;
      regVec_1432 <= 8'h0;
      regVec_1433 <= 8'h0;
      regVec_1434 <= 8'h0;
      regVec_1435 <= 8'h0;
      regVec_1436 <= 8'h0;
      regVec_1437 <= 8'h0;
      regVec_1438 <= 8'h0;
      regVec_1439 <= 8'h0;
      regVec_1440 <= 8'h0;
      regVec_1441 <= 8'h0;
      regVec_1442 <= 8'h0;
      regVec_1443 <= 8'h0;
      regVec_1444 <= 8'h0;
      regVec_1445 <= 8'h0;
      regVec_1446 <= 8'h0;
      regVec_1447 <= 8'h0;
      regVec_1448 <= 8'h0;
      regVec_1449 <= 8'h0;
      regVec_1450 <= 8'h0;
      regVec_1451 <= 8'h0;
      regVec_1452 <= 8'h0;
      regVec_1453 <= 8'h0;
      regVec_1454 <= 8'h0;
      regVec_1455 <= 8'h0;
      regVec_1456 <= 8'h0;
      regVec_1457 <= 8'h0;
      regVec_1458 <= 8'h0;
      regVec_1459 <= 8'h0;
      regVec_1460 <= 8'h0;
      regVec_1461 <= 8'h0;
      regVec_1462 <= 8'h0;
      regVec_1463 <= 8'h0;
      regVec_1464 <= 8'h0;
      regVec_1465 <= 8'h0;
      regVec_1466 <= 8'h0;
      regVec_1467 <= 8'h0;
      regVec_1468 <= 8'h0;
      regVec_1469 <= 8'h0;
      regVec_1470 <= 8'h0;
      regVec_1471 <= 8'h0;
      regVec_1472 <= 8'h0;
      regVec_1473 <= 8'h0;
      regVec_1474 <= 8'h0;
      regVec_1475 <= 8'h0;
      regVec_1476 <= 8'h0;
      regVec_1477 <= 8'h0;
      regVec_1478 <= 8'h0;
      regVec_1479 <= 8'h0;
      regVec_1480 <= 8'h0;
      regVec_1481 <= 8'h0;
      regVec_1482 <= 8'h0;
      regVec_1483 <= 8'h0;
      regVec_1484 <= 8'h0;
      regVec_1485 <= 8'h0;
      regVec_1486 <= 8'h0;
      regVec_1487 <= 8'h0;
      regVec_1488 <= 8'h0;
      regVec_1489 <= 8'h0;
      regVec_1490 <= 8'h0;
      regVec_1491 <= 8'h0;
      regVec_1492 <= 8'h0;
      regVec_1493 <= 8'h0;
      regVec_1494 <= 8'h0;
      regVec_1495 <= 8'h0;
      regVec_1496 <= 8'h0;
      regVec_1497 <= 8'h0;
      regVec_1498 <= 8'h0;
      regVec_1499 <= 8'h0;
      regVec_1500 <= 8'h0;
      regVec_1501 <= 8'h0;
      regVec_1502 <= 8'h0;
      regVec_1503 <= 8'h0;
      regVec_1504 <= 8'h0;
      regVec_1505 <= 8'h0;
      regVec_1506 <= 8'h0;
      regVec_1507 <= 8'h0;
      regVec_1508 <= 8'h0;
      regVec_1509 <= 8'h0;
      regVec_1510 <= 8'h0;
      regVec_1511 <= 8'h0;
      regVec_1512 <= 8'h0;
      regVec_1513 <= 8'h0;
      regVec_1514 <= 8'h0;
      regVec_1515 <= 8'h0;
      regVec_1516 <= 8'h0;
      regVec_1517 <= 8'h0;
      regVec_1518 <= 8'h0;
      regVec_1519 <= 8'h0;
      regVec_1520 <= 8'h0;
      regVec_1521 <= 8'h0;
      regVec_1522 <= 8'h0;
      regVec_1523 <= 8'h0;
      regVec_1524 <= 8'h0;
      regVec_1525 <= 8'h0;
      regVec_1526 <= 8'h0;
      regVec_1527 <= 8'h0;
      regVec_1528 <= 8'h0;
      regVec_1529 <= 8'h0;
      regVec_1530 <= 8'h0;
      regVec_1531 <= 8'h0;
      regVec_1532 <= 8'h0;
      regVec_1533 <= 8'h0;
      regVec_1534 <= 8'h0;
      regVec_1535 <= 8'h0;
      regVec_1536 <= 8'h0;
      regVec_1537 <= 8'h0;
      regVec_1538 <= 8'h0;
      regVec_1539 <= 8'h0;
      regVec_1540 <= 8'h0;
      regVec_1541 <= 8'h0;
      regVec_1542 <= 8'h0;
      regVec_1543 <= 8'h0;
      regVec_1544 <= 8'h0;
      regVec_1545 <= 8'h0;
      regVec_1546 <= 8'h0;
      regVec_1547 <= 8'h0;
      regVec_1548 <= 8'h0;
      regVec_1549 <= 8'h0;
      regVec_1550 <= 8'h0;
      regVec_1551 <= 8'h0;
      regVec_1552 <= 8'h0;
      regVec_1553 <= 8'h0;
      regVec_1554 <= 8'h0;
      regVec_1555 <= 8'h0;
      regVec_1556 <= 8'h0;
      regVec_1557 <= 8'h0;
      regVec_1558 <= 8'h0;
      regVec_1559 <= 8'h0;
      regVec_1560 <= 8'h0;
      regVec_1561 <= 8'h0;
      regVec_1562 <= 8'h0;
      regVec_1563 <= 8'h0;
      regVec_1564 <= 8'h0;
      regVec_1565 <= 8'h0;
      regVec_1566 <= 8'h0;
      regVec_1567 <= 8'h0;
      regVec_1568 <= 8'h0;
      regVec_1569 <= 8'h0;
      regVec_1570 <= 8'h0;
      regVec_1571 <= 8'h0;
      regVec_1572 <= 8'h0;
      regVec_1573 <= 8'h0;
      regVec_1574 <= 8'h0;
      regVec_1575 <= 8'h0;
      regVec_1576 <= 8'h0;
      regVec_1577 <= 8'h0;
      regVec_1578 <= 8'h0;
      regVec_1579 <= 8'h0;
      regVec_1580 <= 8'h0;
      regVec_1581 <= 8'h0;
      regVec_1582 <= 8'h0;
      regVec_1583 <= 8'h0;
      regVec_1584 <= 8'h0;
      regVec_1585 <= 8'h0;
      regVec_1586 <= 8'h0;
      regVec_1587 <= 8'h0;
      regVec_1588 <= 8'h0;
      regVec_1589 <= 8'h0;
      regVec_1590 <= 8'h0;
      regVec_1591 <= 8'h0;
      regVec_1592 <= 8'h0;
      regVec_1593 <= 8'h0;
      regVec_1594 <= 8'h0;
      regVec_1595 <= 8'h0;
      regVec_1596 <= 8'h0;
      regVec_1597 <= 8'h0;
      regVec_1598 <= 8'h0;
      regVec_1599 <= 8'h0;
      regVec_1600 <= 8'h0;
      regVec_1601 <= 8'h0;
      regVec_1602 <= 8'h0;
      regVec_1603 <= 8'h0;
      regVec_1604 <= 8'h0;
      regVec_1605 <= 8'h0;
      regVec_1606 <= 8'h0;
      regVec_1607 <= 8'h0;
      regVec_1608 <= 8'h0;
      regVec_1609 <= 8'h0;
      regVec_1610 <= 8'h0;
      regVec_1611 <= 8'h0;
      regVec_1612 <= 8'h0;
      regVec_1613 <= 8'h0;
      regVec_1614 <= 8'h0;
      regVec_1615 <= 8'h0;
      regVec_1616 <= 8'h0;
      regVec_1617 <= 8'h0;
      regVec_1618 <= 8'h0;
      regVec_1619 <= 8'h0;
      regVec_1620 <= 8'h0;
      regVec_1621 <= 8'h0;
      regVec_1622 <= 8'h0;
      regVec_1623 <= 8'h0;
      regVec_1624 <= 8'h0;
      regVec_1625 <= 8'h0;
      regVec_1626 <= 8'h0;
      regVec_1627 <= 8'h0;
      regVec_1628 <= 8'h0;
      regVec_1629 <= 8'h0;
      regVec_1630 <= 8'h0;
      regVec_1631 <= 8'h0;
      regVec_1632 <= 8'h0;
      regVec_1633 <= 8'h0;
      regVec_1634 <= 8'h0;
      regVec_1635 <= 8'h0;
      regVec_1636 <= 8'h0;
      regVec_1637 <= 8'h0;
      regVec_1638 <= 8'h0;
      regVec_1639 <= 8'h0;
      regVec_1640 <= 8'h0;
      regVec_1641 <= 8'h0;
      regVec_1642 <= 8'h0;
      regVec_1643 <= 8'h0;
      regVec_1644 <= 8'h0;
      regVec_1645 <= 8'h0;
      regVec_1646 <= 8'h0;
      regVec_1647 <= 8'h0;
      regVec_1648 <= 8'h0;
      regVec_1649 <= 8'h0;
      regVec_1650 <= 8'h0;
      regVec_1651 <= 8'h0;
      regVec_1652 <= 8'h0;
      regVec_1653 <= 8'h0;
      regVec_1654 <= 8'h0;
      regVec_1655 <= 8'h0;
      regVec_1656 <= 8'h0;
      regVec_1657 <= 8'h0;
      regVec_1658 <= 8'h0;
      regVec_1659 <= 8'h0;
      regVec_1660 <= 8'h0;
      regVec_1661 <= 8'h0;
      regVec_1662 <= 8'h0;
      regVec_1663 <= 8'h0;
      regVec_1664 <= 8'h0;
      regVec_1665 <= 8'h0;
      regVec_1666 <= 8'h0;
      regVec_1667 <= 8'h0;
      regVec_1668 <= 8'h0;
      regVec_1669 <= 8'h0;
      regVec_1670 <= 8'h0;
      regVec_1671 <= 8'h0;
      regVec_1672 <= 8'h0;
      regVec_1673 <= 8'h0;
      regVec_1674 <= 8'h0;
      regVec_1675 <= 8'h0;
      regVec_1676 <= 8'h0;
      regVec_1677 <= 8'h0;
      regVec_1678 <= 8'h0;
      regVec_1679 <= 8'h0;
      regVec_1680 <= 8'h0;
      regVec_1681 <= 8'h0;
      regVec_1682 <= 8'h0;
      regVec_1683 <= 8'h0;
      regVec_1684 <= 8'h0;
      regVec_1685 <= 8'h0;
      regVec_1686 <= 8'h0;
      regVec_1687 <= 8'h0;
      regVec_1688 <= 8'h0;
      regVec_1689 <= 8'h0;
      regVec_1690 <= 8'h0;
      regVec_1691 <= 8'h0;
      regVec_1692 <= 8'h0;
      regVec_1693 <= 8'h0;
      regVec_1694 <= 8'h0;
      regVec_1695 <= 8'h0;
      regVec_1696 <= 8'h0;
      regVec_1697 <= 8'h0;
      regVec_1698 <= 8'h0;
      regVec_1699 <= 8'h0;
      regVec_1700 <= 8'h0;
      regVec_1701 <= 8'h0;
      regVec_1702 <= 8'h0;
      regVec_1703 <= 8'h0;
      regVec_1704 <= 8'h0;
      regVec_1705 <= 8'h0;
      regVec_1706 <= 8'h0;
      regVec_1707 <= 8'h0;
      regVec_1708 <= 8'h0;
      regVec_1709 <= 8'h0;
      regVec_1710 <= 8'h0;
      regVec_1711 <= 8'h0;
      regVec_1712 <= 8'h0;
      regVec_1713 <= 8'h0;
      regVec_1714 <= 8'h0;
      regVec_1715 <= 8'h0;
      regVec_1716 <= 8'h0;
      regVec_1717 <= 8'h0;
      regVec_1718 <= 8'h0;
      regVec_1719 <= 8'h0;
      regVec_1720 <= 8'h0;
      regVec_1721 <= 8'h0;
      regVec_1722 <= 8'h0;
      regVec_1723 <= 8'h0;
      regVec_1724 <= 8'h0;
      regVec_1725 <= 8'h0;
      regVec_1726 <= 8'h0;
      regVec_1727 <= 8'h0;
      regVec_1728 <= 8'h0;
      regVec_1729 <= 8'h0;
      regVec_1730 <= 8'h0;
      regVec_1731 <= 8'h0;
      regVec_1732 <= 8'h0;
      regVec_1733 <= 8'h0;
      regVec_1734 <= 8'h0;
      regVec_1735 <= 8'h0;
      regVec_1736 <= 8'h0;
      regVec_1737 <= 8'h0;
      regVec_1738 <= 8'h0;
      regVec_1739 <= 8'h0;
      regVec_1740 <= 8'h0;
      regVec_1741 <= 8'h0;
      regVec_1742 <= 8'h0;
      regVec_1743 <= 8'h0;
      regVec_1744 <= 8'h0;
      regVec_1745 <= 8'h0;
      regVec_1746 <= 8'h0;
      regVec_1747 <= 8'h0;
      regVec_1748 <= 8'h0;
      regVec_1749 <= 8'h0;
      regVec_1750 <= 8'h0;
      regVec_1751 <= 8'h0;
      regVec_1752 <= 8'h0;
      regVec_1753 <= 8'h0;
      regVec_1754 <= 8'h0;
      regVec_1755 <= 8'h0;
      regVec_1756 <= 8'h0;
      regVec_1757 <= 8'h0;
      regVec_1758 <= 8'h0;
      regVec_1759 <= 8'h0;
      regVec_1760 <= 8'h0;
      regVec_1761 <= 8'h0;
      regVec_1762 <= 8'h0;
      regVec_1763 <= 8'h0;
      regVec_1764 <= 8'h0;
      regVec_1765 <= 8'h0;
      regVec_1766 <= 8'h0;
      regVec_1767 <= 8'h0;
      regVec_1768 <= 8'h0;
      regVec_1769 <= 8'h0;
      regVec_1770 <= 8'h0;
      regVec_1771 <= 8'h0;
      regVec_1772 <= 8'h0;
      regVec_1773 <= 8'h0;
      regVec_1774 <= 8'h0;
      regVec_1775 <= 8'h0;
      regVec_1776 <= 8'h0;
      regVec_1777 <= 8'h0;
      regVec_1778 <= 8'h0;
      regVec_1779 <= 8'h0;
      regVec_1780 <= 8'h0;
      regVec_1781 <= 8'h0;
      regVec_1782 <= 8'h0;
      regVec_1783 <= 8'h0;
      regVec_1784 <= 8'h0;
      regVec_1785 <= 8'h0;
      regVec_1786 <= 8'h0;
      regVec_1787 <= 8'h0;
      regVec_1788 <= 8'h0;
      regVec_1789 <= 8'h0;
      regVec_1790 <= 8'h0;
      regVec_1791 <= 8'h0;
      regVec_1792 <= 8'h0;
      regVec_1793 <= 8'h0;
      regVec_1794 <= 8'h0;
      regVec_1795 <= 8'h0;
      regVec_1796 <= 8'h0;
      regVec_1797 <= 8'h0;
      regVec_1798 <= 8'h0;
      regVec_1799 <= 8'h0;
      regVec_1800 <= 8'h0;
      regVec_1801 <= 8'h0;
      regVec_1802 <= 8'h0;
      regVec_1803 <= 8'h0;
      regVec_1804 <= 8'h0;
      regVec_1805 <= 8'h0;
      regVec_1806 <= 8'h0;
      regVec_1807 <= 8'h0;
      regVec_1808 <= 8'h0;
      regVec_1809 <= 8'h0;
      regVec_1810 <= 8'h0;
      regVec_1811 <= 8'h0;
      regVec_1812 <= 8'h0;
      regVec_1813 <= 8'h0;
      regVec_1814 <= 8'h0;
      regVec_1815 <= 8'h0;
      regVec_1816 <= 8'h0;
      regVec_1817 <= 8'h0;
      regVec_1818 <= 8'h0;
      regVec_1819 <= 8'h0;
      regVec_1820 <= 8'h0;
      regVec_1821 <= 8'h0;
      regVec_1822 <= 8'h0;
      regVec_1823 <= 8'h0;
      regVec_1824 <= 8'h0;
      regVec_1825 <= 8'h0;
      regVec_1826 <= 8'h0;
      regVec_1827 <= 8'h0;
      regVec_1828 <= 8'h0;
      regVec_1829 <= 8'h0;
      regVec_1830 <= 8'h0;
      regVec_1831 <= 8'h0;
      regVec_1832 <= 8'h0;
      regVec_1833 <= 8'h0;
      regVec_1834 <= 8'h0;
      regVec_1835 <= 8'h0;
      regVec_1836 <= 8'h0;
      regVec_1837 <= 8'h0;
      regVec_1838 <= 8'h0;
      regVec_1839 <= 8'h0;
      regVec_1840 <= 8'h0;
      regVec_1841 <= 8'h0;
      regVec_1842 <= 8'h0;
      regVec_1843 <= 8'h0;
      regVec_1844 <= 8'h0;
      regVec_1845 <= 8'h0;
      regVec_1846 <= 8'h0;
      regVec_1847 <= 8'h0;
      regVec_1848 <= 8'h0;
      regVec_1849 <= 8'h0;
      regVec_1850 <= 8'h0;
      regVec_1851 <= 8'h0;
      regVec_1852 <= 8'h0;
      regVec_1853 <= 8'h0;
      regVec_1854 <= 8'h0;
      regVec_1855 <= 8'h0;
      regVec_1856 <= 8'h0;
      regVec_1857 <= 8'h0;
      regVec_1858 <= 8'h0;
      regVec_1859 <= 8'h0;
      regVec_1860 <= 8'h0;
      regVec_1861 <= 8'h0;
      regVec_1862 <= 8'h0;
      regVec_1863 <= 8'h0;
      regVec_1864 <= 8'h0;
      regVec_1865 <= 8'h0;
      regVec_1866 <= 8'h0;
      regVec_1867 <= 8'h0;
      regVec_1868 <= 8'h0;
      regVec_1869 <= 8'h0;
      regVec_1870 <= 8'h0;
      regVec_1871 <= 8'h0;
      regVec_1872 <= 8'h0;
      regVec_1873 <= 8'h0;
      regVec_1874 <= 8'h0;
      regVec_1875 <= 8'h0;
      regVec_1876 <= 8'h0;
      regVec_1877 <= 8'h0;
      regVec_1878 <= 8'h0;
      regVec_1879 <= 8'h0;
      regVec_1880 <= 8'h0;
      regVec_1881 <= 8'h0;
      regVec_1882 <= 8'h0;
      regVec_1883 <= 8'h0;
      regVec_1884 <= 8'h0;
      regVec_1885 <= 8'h0;
      regVec_1886 <= 8'h0;
      regVec_1887 <= 8'h0;
      regVec_1888 <= 8'h0;
      regVec_1889 <= 8'h0;
      regVec_1890 <= 8'h0;
      regVec_1891 <= 8'h0;
      regVec_1892 <= 8'h0;
      regVec_1893 <= 8'h0;
      regVec_1894 <= 8'h0;
      regVec_1895 <= 8'h0;
      regVec_1896 <= 8'h0;
      regVec_1897 <= 8'h0;
      regVec_1898 <= 8'h0;
      regVec_1899 <= 8'h0;
      regVec_1900 <= 8'h0;
      regVec_1901 <= 8'h0;
      regVec_1902 <= 8'h0;
      regVec_1903 <= 8'h0;
      regVec_1904 <= 8'h0;
      regVec_1905 <= 8'h0;
      regVec_1906 <= 8'h0;
      regVec_1907 <= 8'h0;
      regVec_1908 <= 8'h0;
      regVec_1909 <= 8'h0;
      regVec_1910 <= 8'h0;
      regVec_1911 <= 8'h0;
      regVec_1912 <= 8'h0;
      regVec_1913 <= 8'h0;
      regVec_1914 <= 8'h0;
      regVec_1915 <= 8'h0;
      regVec_1916 <= 8'h0;
      regVec_1917 <= 8'h0;
      regVec_1918 <= 8'h0;
      regVec_1919 <= 8'h0;
      regVec_1920 <= 8'h0;
      regVec_1921 <= 8'h0;
      regVec_1922 <= 8'h0;
      regVec_1923 <= 8'h0;
      regVec_1924 <= 8'h0;
      regVec_1925 <= 8'h0;
      regVec_1926 <= 8'h0;
      regVec_1927 <= 8'h0;
      regVec_1928 <= 8'h0;
      regVec_1929 <= 8'h0;
      regVec_1930 <= 8'h0;
      regVec_1931 <= 8'h0;
      regVec_1932 <= 8'h0;
      regVec_1933 <= 8'h0;
      regVec_1934 <= 8'h0;
      regVec_1935 <= 8'h0;
      regVec_1936 <= 8'h0;
      regVec_1937 <= 8'h0;
      regVec_1938 <= 8'h0;
      regVec_1939 <= 8'h0;
      regVec_1940 <= 8'h0;
      regVec_1941 <= 8'h0;
      regVec_1942 <= 8'h0;
      regVec_1943 <= 8'h0;
      regVec_1944 <= 8'h0;
      regVec_1945 <= 8'h0;
      regVec_1946 <= 8'h0;
      regVec_1947 <= 8'h0;
      regVec_1948 <= 8'h0;
      regVec_1949 <= 8'h0;
      regVec_1950 <= 8'h0;
      regVec_1951 <= 8'h0;
      regVec_1952 <= 8'h0;
      regVec_1953 <= 8'h0;
      regVec_1954 <= 8'h0;
      regVec_1955 <= 8'h0;
      regVec_1956 <= 8'h0;
      regVec_1957 <= 8'h0;
      regVec_1958 <= 8'h0;
      regVec_1959 <= 8'h0;
      regVec_1960 <= 8'h0;
      regVec_1961 <= 8'h0;
      regVec_1962 <= 8'h0;
      regVec_1963 <= 8'h0;
      regVec_1964 <= 8'h0;
      regVec_1965 <= 8'h0;
      regVec_1966 <= 8'h0;
      regVec_1967 <= 8'h0;
      regVec_1968 <= 8'h0;
      regVec_1969 <= 8'h0;
      regVec_1970 <= 8'h0;
      regVec_1971 <= 8'h0;
      regVec_1972 <= 8'h0;
      regVec_1973 <= 8'h0;
      regVec_1974 <= 8'h0;
      regVec_1975 <= 8'h0;
      regVec_1976 <= 8'h0;
      regVec_1977 <= 8'h0;
      regVec_1978 <= 8'h0;
      regVec_1979 <= 8'h0;
      regVec_1980 <= 8'h0;
      regVec_1981 <= 8'h0;
      regVec_1982 <= 8'h0;
      regVec_1983 <= 8'h0;
      regVec_1984 <= 8'h0;
      regVec_1985 <= 8'h0;
      regVec_1986 <= 8'h0;
      regVec_1987 <= 8'h0;
      regVec_1988 <= 8'h0;
      regVec_1989 <= 8'h0;
      regVec_1990 <= 8'h0;
      regVec_1991 <= 8'h0;
      regVec_1992 <= 8'h0;
      regVec_1993 <= 8'h0;
      regVec_1994 <= 8'h0;
      regVec_1995 <= 8'h0;
      regVec_1996 <= 8'h0;
      regVec_1997 <= 8'h0;
      regVec_1998 <= 8'h0;
      regVec_1999 <= 8'h0;
      regVec_2000 <= 8'h0;
      regVec_2001 <= 8'h0;
      regVec_2002 <= 8'h0;
      regVec_2003 <= 8'h0;
      regVec_2004 <= 8'h0;
      regVec_2005 <= 8'h0;
      regVec_2006 <= 8'h0;
      regVec_2007 <= 8'h0;
      regVec_2008 <= 8'h0;
      regVec_2009 <= 8'h0;
      regVec_2010 <= 8'h0;
      regVec_2011 <= 8'h0;
      regVec_2012 <= 8'h0;
      regVec_2013 <= 8'h0;
      regVec_2014 <= 8'h0;
      regVec_2015 <= 8'h0;
      regVec_2016 <= 8'h0;
      regVec_2017 <= 8'h0;
      regVec_2018 <= 8'h0;
      regVec_2019 <= 8'h0;
      regVec_2020 <= 8'h0;
      regVec_2021 <= 8'h0;
      regVec_2022 <= 8'h0;
      regVec_2023 <= 8'h0;
      regVec_2024 <= 8'h0;
      regVec_2025 <= 8'h0;
      regVec_2026 <= 8'h0;
      regVec_2027 <= 8'h0;
      regVec_2028 <= 8'h0;
      regVec_2029 <= 8'h0;
      regVec_2030 <= 8'h0;
      regVec_2031 <= 8'h0;
      regVec_2032 <= 8'h0;
      regVec_2033 <= 8'h0;
      regVec_2034 <= 8'h0;
      regVec_2035 <= 8'h0;
      regVec_2036 <= 8'h0;
      regVec_2037 <= 8'h0;
      regVec_2038 <= 8'h0;
      regVec_2039 <= 8'h0;
      regVec_2040 <= 8'h0;
      regVec_2041 <= 8'h0;
      regVec_2042 <= 8'h0;
      regVec_2043 <= 8'h0;
      regVec_2044 <= 8'h0;
      regVec_2045 <= 8'h0;
      regVec_2046 <= 8'h0;
      regVec_2047 <= 8'h0;
      regVec_2048 <= 8'h0;
      regVec_2049 <= 8'h0;
      regVec_2050 <= 8'h0;
      regVec_2051 <= 8'h0;
      regVec_2052 <= 8'h0;
      regVec_2053 <= 8'h0;
      regVec_2054 <= 8'h0;
      regVec_2055 <= 8'h0;
      regVec_2056 <= 8'h0;
      regVec_2057 <= 8'h0;
      regVec_2058 <= 8'h0;
      regVec_2059 <= 8'h0;
      regVec_2060 <= 8'h0;
      regVec_2061 <= 8'h0;
      regVec_2062 <= 8'h0;
      regVec_2063 <= 8'h0;
      regVec_2064 <= 8'h0;
      regVec_2065 <= 8'h0;
      regVec_2066 <= 8'h0;
      regVec_2067 <= 8'h0;
      regVec_2068 <= 8'h0;
      regVec_2069 <= 8'h0;
      regVec_2070 <= 8'h0;
      regVec_2071 <= 8'h0;
      regVec_2072 <= 8'h0;
      regVec_2073 <= 8'h0;
      regVec_2074 <= 8'h0;
      regVec_2075 <= 8'h0;
      regVec_2076 <= 8'h0;
      regVec_2077 <= 8'h0;
      regVec_2078 <= 8'h0;
      regVec_2079 <= 8'h0;
      regVec_2080 <= 8'h0;
      regVec_2081 <= 8'h0;
      regVec_2082 <= 8'h0;
      regVec_2083 <= 8'h0;
      regVec_2084 <= 8'h0;
      regVec_2085 <= 8'h0;
      regVec_2086 <= 8'h0;
      regVec_2087 <= 8'h0;
      regVec_2088 <= 8'h0;
      regVec_2089 <= 8'h0;
      regVec_2090 <= 8'h0;
      regVec_2091 <= 8'h0;
      regVec_2092 <= 8'h0;
      regVec_2093 <= 8'h0;
      regVec_2094 <= 8'h0;
      regVec_2095 <= 8'h0;
      regVec_2096 <= 8'h0;
      regVec_2097 <= 8'h0;
      regVec_2098 <= 8'h0;
      regVec_2099 <= 8'h0;
      regVec_2100 <= 8'h0;
      regVec_2101 <= 8'h0;
      regVec_2102 <= 8'h0;
      regVec_2103 <= 8'h0;
      regVec_2104 <= 8'h0;
      regVec_2105 <= 8'h0;
      regVec_2106 <= 8'h0;
      regVec_2107 <= 8'h0;
      regVec_2108 <= 8'h0;
      regVec_2109 <= 8'h0;
      regVec_2110 <= 8'h0;
      regVec_2111 <= 8'h0;
      regVec_2112 <= 8'h0;
      regVec_2113 <= 8'h0;
      regVec_2114 <= 8'h0;
      regVec_2115 <= 8'h0;
      regVec_2116 <= 8'h0;
      regVec_2117 <= 8'h0;
      regVec_2118 <= 8'h0;
      regVec_2119 <= 8'h0;
      regVec_2120 <= 8'h0;
      regVec_2121 <= 8'h0;
      regVec_2122 <= 8'h0;
      regVec_2123 <= 8'h0;
      regVec_2124 <= 8'h0;
      regVec_2125 <= 8'h0;
      regVec_2126 <= 8'h0;
      regVec_2127 <= 8'h0;
      regVec_2128 <= 8'h0;
      regVec_2129 <= 8'h0;
      regVec_2130 <= 8'h0;
      regVec_2131 <= 8'h0;
      regVec_2132 <= 8'h0;
      regVec_2133 <= 8'h0;
      regVec_2134 <= 8'h0;
      regVec_2135 <= 8'h0;
      regVec_2136 <= 8'h0;
      regVec_2137 <= 8'h0;
      regVec_2138 <= 8'h0;
      regVec_2139 <= 8'h0;
      regVec_2140 <= 8'h0;
      regVec_2141 <= 8'h0;
      regVec_2142 <= 8'h0;
      regVec_2143 <= 8'h0;
      regVec_2144 <= 8'h0;
      regVec_2145 <= 8'h0;
      regVec_2146 <= 8'h0;
      regVec_2147 <= 8'h0;
      regVec_2148 <= 8'h0;
      regVec_2149 <= 8'h0;
      regVec_2150 <= 8'h0;
      regVec_2151 <= 8'h0;
      regVec_2152 <= 8'h0;
      regVec_2153 <= 8'h0;
      regVec_2154 <= 8'h0;
      regVec_2155 <= 8'h0;
      regVec_2156 <= 8'h0;
      regVec_2157 <= 8'h0;
      regVec_2158 <= 8'h0;
      regVec_2159 <= 8'h0;
      regVec_2160 <= 8'h0;
      regVec_2161 <= 8'h0;
      regVec_2162 <= 8'h0;
      regVec_2163 <= 8'h0;
      regVec_2164 <= 8'h0;
      regVec_2165 <= 8'h0;
      regVec_2166 <= 8'h0;
      regVec_2167 <= 8'h0;
      regVec_2168 <= 8'h0;
      regVec_2169 <= 8'h0;
      regVec_2170 <= 8'h0;
      regVec_2171 <= 8'h0;
      regVec_2172 <= 8'h0;
      regVec_2173 <= 8'h0;
      regVec_2174 <= 8'h0;
      regVec_2175 <= 8'h0;
      regVec_2176 <= 8'h0;
      regVec_2177 <= 8'h0;
      regVec_2178 <= 8'h0;
      regVec_2179 <= 8'h0;
      regVec_2180 <= 8'h0;
      regVec_2181 <= 8'h0;
      regVec_2182 <= 8'h0;
      regVec_2183 <= 8'h0;
      regVec_2184 <= 8'h0;
      regVec_2185 <= 8'h0;
      regVec_2186 <= 8'h0;
      regVec_2187 <= 8'h0;
      regVec_2188 <= 8'h0;
      regVec_2189 <= 8'h0;
      regVec_2190 <= 8'h0;
      regVec_2191 <= 8'h0;
      regVec_2192 <= 8'h0;
      regVec_2193 <= 8'h0;
      regVec_2194 <= 8'h0;
      regVec_2195 <= 8'h0;
      regVec_2196 <= 8'h0;
      regVec_2197 <= 8'h0;
      regVec_2198 <= 8'h0;
      regVec_2199 <= 8'h0;
      regVec_2200 <= 8'h0;
      regVec_2201 <= 8'h0;
      regVec_2202 <= 8'h0;
      regVec_2203 <= 8'h0;
      regVec_2204 <= 8'h0;
      regVec_2205 <= 8'h0;
      regVec_2206 <= 8'h0;
      regVec_2207 <= 8'h0;
      regVec_2208 <= 8'h0;
      regVec_2209 <= 8'h0;
      regVec_2210 <= 8'h0;
      regVec_2211 <= 8'h0;
      regVec_2212 <= 8'h0;
      regVec_2213 <= 8'h0;
      regVec_2214 <= 8'h0;
      regVec_2215 <= 8'h0;
      regVec_2216 <= 8'h0;
      regVec_2217 <= 8'h0;
      regVec_2218 <= 8'h0;
      regVec_2219 <= 8'h0;
      regVec_2220 <= 8'h0;
      regVec_2221 <= 8'h0;
      regVec_2222 <= 8'h0;
      regVec_2223 <= 8'h0;
      regVec_2224 <= 8'h0;
      regVec_2225 <= 8'h0;
      regVec_2226 <= 8'h0;
      regVec_2227 <= 8'h0;
      regVec_2228 <= 8'h0;
      regVec_2229 <= 8'h0;
      regVec_2230 <= 8'h0;
      regVec_2231 <= 8'h0;
      regVec_2232 <= 8'h0;
      regVec_2233 <= 8'h0;
      regVec_2234 <= 8'h0;
      regVec_2235 <= 8'h0;
      regVec_2236 <= 8'h0;
      regVec_2237 <= 8'h0;
      regVec_2238 <= 8'h0;
      regVec_2239 <= 8'h0;
      regVec_2240 <= 8'h0;
      regVec_2241 <= 8'h0;
      regVec_2242 <= 8'h0;
      regVec_2243 <= 8'h0;
      regVec_2244 <= 8'h0;
      regVec_2245 <= 8'h0;
      regVec_2246 <= 8'h0;
      regVec_2247 <= 8'h0;
      regVec_2248 <= 8'h0;
      regVec_2249 <= 8'h0;
      regVec_2250 <= 8'h0;
      regVec_2251 <= 8'h0;
      regVec_2252 <= 8'h0;
      regVec_2253 <= 8'h0;
      regVec_2254 <= 8'h0;
      regVec_2255 <= 8'h0;
      regVec_2256 <= 8'h0;
      regVec_2257 <= 8'h0;
      regVec_2258 <= 8'h0;
      regVec_2259 <= 8'h0;
      regVec_2260 <= 8'h0;
      regVec_2261 <= 8'h0;
      regVec_2262 <= 8'h0;
      regVec_2263 <= 8'h0;
      regVec_2264 <= 8'h0;
      regVec_2265 <= 8'h0;
      regVec_2266 <= 8'h0;
      regVec_2267 <= 8'h0;
      regVec_2268 <= 8'h0;
      regVec_2269 <= 8'h0;
      regVec_2270 <= 8'h0;
      regVec_2271 <= 8'h0;
      regVec_2272 <= 8'h0;
      regVec_2273 <= 8'h0;
      regVec_2274 <= 8'h0;
      regVec_2275 <= 8'h0;
      regVec_2276 <= 8'h0;
      regVec_2277 <= 8'h0;
      regVec_2278 <= 8'h0;
      regVec_2279 <= 8'h0;
      regVec_2280 <= 8'h0;
      regVec_2281 <= 8'h0;
      regVec_2282 <= 8'h0;
      regVec_2283 <= 8'h0;
      regVec_2284 <= 8'h0;
      regVec_2285 <= 8'h0;
      regVec_2286 <= 8'h0;
      regVec_2287 <= 8'h0;
      regVec_2288 <= 8'h0;
      regVec_2289 <= 8'h0;
      regVec_2290 <= 8'h0;
      regVec_2291 <= 8'h0;
      regVec_2292 <= 8'h0;
      regVec_2293 <= 8'h0;
      regVec_2294 <= 8'h0;
      regVec_2295 <= 8'h0;
      regVec_2296 <= 8'h0;
      regVec_2297 <= 8'h0;
      regVec_2298 <= 8'h0;
      regVec_2299 <= 8'h0;
      regVec_2300 <= 8'h0;
      regVec_2301 <= 8'h0;
      regVec_2302 <= 8'h0;
      regVec_2303 <= 8'h0;
      regVec_2304 <= 8'h0;
      regVec_2305 <= 8'h0;
      regVec_2306 <= 8'h0;
      regVec_2307 <= 8'h0;
      regVec_2308 <= 8'h0;
      regVec_2309 <= 8'h0;
      regVec_2310 <= 8'h0;
      regVec_2311 <= 8'h0;
      regVec_2312 <= 8'h0;
      regVec_2313 <= 8'h0;
      regVec_2314 <= 8'h0;
      regVec_2315 <= 8'h0;
      regVec_2316 <= 8'h0;
      regVec_2317 <= 8'h0;
      regVec_2318 <= 8'h0;
      regVec_2319 <= 8'h0;
      regVec_2320 <= 8'h0;
      regVec_2321 <= 8'h0;
      regVec_2322 <= 8'h0;
      regVec_2323 <= 8'h0;
      regVec_2324 <= 8'h0;
      regVec_2325 <= 8'h0;
      regVec_2326 <= 8'h0;
      regVec_2327 <= 8'h0;
      regVec_2328 <= 8'h0;
      regVec_2329 <= 8'h0;
      regVec_2330 <= 8'h0;
      regVec_2331 <= 8'h0;
      regVec_2332 <= 8'h0;
      regVec_2333 <= 8'h0;
      regVec_2334 <= 8'h0;
      regVec_2335 <= 8'h0;
      regVec_2336 <= 8'h0;
      regVec_2337 <= 8'h0;
      regVec_2338 <= 8'h0;
      regVec_2339 <= 8'h0;
      regVec_2340 <= 8'h0;
      regVec_2341 <= 8'h0;
      regVec_2342 <= 8'h0;
      regVec_2343 <= 8'h0;
      regVec_2344 <= 8'h0;
      regVec_2345 <= 8'h0;
      regVec_2346 <= 8'h0;
      regVec_2347 <= 8'h0;
      regVec_2348 <= 8'h0;
      regVec_2349 <= 8'h0;
      regVec_2350 <= 8'h0;
      regVec_2351 <= 8'h0;
      regVec_2352 <= 8'h0;
      regVec_2353 <= 8'h0;
      regVec_2354 <= 8'h0;
      regVec_2355 <= 8'h0;
      regVec_2356 <= 8'h0;
      regVec_2357 <= 8'h0;
      regVec_2358 <= 8'h0;
      regVec_2359 <= 8'h0;
      regVec_2360 <= 8'h0;
      regVec_2361 <= 8'h0;
      regVec_2362 <= 8'h0;
      regVec_2363 <= 8'h0;
      regVec_2364 <= 8'h0;
      regVec_2365 <= 8'h0;
      regVec_2366 <= 8'h0;
      regVec_2367 <= 8'h0;
      regVec_2368 <= 8'h0;
      regVec_2369 <= 8'h0;
      regVec_2370 <= 8'h0;
      regVec_2371 <= 8'h0;
      regVec_2372 <= 8'h0;
      regVec_2373 <= 8'h0;
      regVec_2374 <= 8'h0;
      regVec_2375 <= 8'h0;
      regVec_2376 <= 8'h0;
      regVec_2377 <= 8'h0;
      regVec_2378 <= 8'h0;
      regVec_2379 <= 8'h0;
      regVec_2380 <= 8'h0;
      regVec_2381 <= 8'h0;
      regVec_2382 <= 8'h0;
      regVec_2383 <= 8'h0;
      regVec_2384 <= 8'h0;
      regVec_2385 <= 8'h0;
      regVec_2386 <= 8'h0;
      regVec_2387 <= 8'h0;
      regVec_2388 <= 8'h0;
      regVec_2389 <= 8'h0;
      regVec_2390 <= 8'h0;
      regVec_2391 <= 8'h0;
      regVec_2392 <= 8'h0;
      regVec_2393 <= 8'h0;
      regVec_2394 <= 8'h0;
      regVec_2395 <= 8'h0;
      regVec_2396 <= 8'h0;
      regVec_2397 <= 8'h0;
      regVec_2398 <= 8'h0;
      regVec_2399 <= 8'h0;
      regVec_2400 <= 8'h0;
      regVec_2401 <= 8'h0;
      regVec_2402 <= 8'h0;
      regVec_2403 <= 8'h0;
      regVec_2404 <= 8'h0;
      regVec_2405 <= 8'h0;
      regVec_2406 <= 8'h0;
      regVec_2407 <= 8'h0;
      regVec_2408 <= 8'h0;
      regVec_2409 <= 8'h0;
      regVec_2410 <= 8'h0;
      regVec_2411 <= 8'h0;
      regVec_2412 <= 8'h0;
      regVec_2413 <= 8'h0;
      regVec_2414 <= 8'h0;
      regVec_2415 <= 8'h0;
      regVec_2416 <= 8'h0;
      regVec_2417 <= 8'h0;
      regVec_2418 <= 8'h0;
      regVec_2419 <= 8'h0;
      regVec_2420 <= 8'h0;
      regVec_2421 <= 8'h0;
      regVec_2422 <= 8'h0;
      regVec_2423 <= 8'h0;
      regVec_2424 <= 8'h0;
      regVec_2425 <= 8'h0;
      regVec_2426 <= 8'h0;
      regVec_2427 <= 8'h0;
      regVec_2428 <= 8'h0;
      regVec_2429 <= 8'h0;
      regVec_2430 <= 8'h0;
      regVec_2431 <= 8'h0;
      regVec_2432 <= 8'h0;
      regVec_2433 <= 8'h0;
      regVec_2434 <= 8'h0;
      regVec_2435 <= 8'h0;
      regVec_2436 <= 8'h0;
      regVec_2437 <= 8'h0;
      regVec_2438 <= 8'h0;
      regVec_2439 <= 8'h0;
      regVec_2440 <= 8'h0;
      regVec_2441 <= 8'h0;
      regVec_2442 <= 8'h0;
      regVec_2443 <= 8'h0;
      regVec_2444 <= 8'h0;
      regVec_2445 <= 8'h0;
      regVec_2446 <= 8'h0;
      regVec_2447 <= 8'h0;
      regVec_2448 <= 8'h0;
      regVec_2449 <= 8'h0;
      regVec_2450 <= 8'h0;
      regVec_2451 <= 8'h0;
      regVec_2452 <= 8'h0;
      regVec_2453 <= 8'h0;
      regVec_2454 <= 8'h0;
      regVec_2455 <= 8'h0;
      regVec_2456 <= 8'h0;
      regVec_2457 <= 8'h0;
      regVec_2458 <= 8'h0;
      regVec_2459 <= 8'h0;
      regVec_2460 <= 8'h0;
      regVec_2461 <= 8'h0;
      regVec_2462 <= 8'h0;
      regVec_2463 <= 8'h0;
      regVec_2464 <= 8'h0;
      regVec_2465 <= 8'h0;
      regVec_2466 <= 8'h0;
      regVec_2467 <= 8'h0;
      regVec_2468 <= 8'h0;
      regVec_2469 <= 8'h0;
      regVec_2470 <= 8'h0;
      regVec_2471 <= 8'h0;
      regVec_2472 <= 8'h0;
      regVec_2473 <= 8'h0;
      regVec_2474 <= 8'h0;
      regVec_2475 <= 8'h0;
      regVec_2476 <= 8'h0;
      regVec_2477 <= 8'h0;
      regVec_2478 <= 8'h0;
      regVec_2479 <= 8'h0;
      regVec_2480 <= 8'h0;
      regVec_2481 <= 8'h0;
      regVec_2482 <= 8'h0;
      regVec_2483 <= 8'h0;
      regVec_2484 <= 8'h0;
      regVec_2485 <= 8'h0;
      regVec_2486 <= 8'h0;
      regVec_2487 <= 8'h0;
      regVec_2488 <= 8'h0;
      regVec_2489 <= 8'h0;
      regVec_2490 <= 8'h0;
      regVec_2491 <= 8'h0;
      regVec_2492 <= 8'h0;
      regVec_2493 <= 8'h0;
      regVec_2494 <= 8'h0;
      regVec_2495 <= 8'h0;
      regVec_2496 <= 8'h0;
      regVec_2497 <= 8'h0;
      regVec_2498 <= 8'h0;
      regVec_2499 <= 8'h0;
      regVec_2500 <= 8'h0;
      regVec_2501 <= 8'h0;
      regVec_2502 <= 8'h0;
      regVec_2503 <= 8'h0;
      regVec_2504 <= 8'h0;
      regVec_2505 <= 8'h0;
      regVec_2506 <= 8'h0;
      regVec_2507 <= 8'h0;
      regVec_2508 <= 8'h0;
      regVec_2509 <= 8'h0;
      regVec_2510 <= 8'h0;
      regVec_2511 <= 8'h0;
      regVec_2512 <= 8'h0;
      regVec_2513 <= 8'h0;
      regVec_2514 <= 8'h0;
      regVec_2515 <= 8'h0;
      regVec_2516 <= 8'h0;
      regVec_2517 <= 8'h0;
      regVec_2518 <= 8'h0;
      regVec_2519 <= 8'h0;
      regVec_2520 <= 8'h0;
      regVec_2521 <= 8'h0;
      regVec_2522 <= 8'h0;
      regVec_2523 <= 8'h0;
      regVec_2524 <= 8'h0;
      regVec_2525 <= 8'h0;
      regVec_2526 <= 8'h0;
      regVec_2527 <= 8'h0;
      regVec_2528 <= 8'h0;
      regVec_2529 <= 8'h0;
      regVec_2530 <= 8'h0;
      regVec_2531 <= 8'h0;
      regVec_2532 <= 8'h0;
      regVec_2533 <= 8'h0;
      regVec_2534 <= 8'h0;
      regVec_2535 <= 8'h0;
      regVec_2536 <= 8'h0;
      regVec_2537 <= 8'h0;
      regVec_2538 <= 8'h0;
      regVec_2539 <= 8'h0;
      regVec_2540 <= 8'h0;
      regVec_2541 <= 8'h0;
      regVec_2542 <= 8'h0;
      regVec_2543 <= 8'h0;
      regVec_2544 <= 8'h0;
      regVec_2545 <= 8'h0;
      regVec_2546 <= 8'h0;
      regVec_2547 <= 8'h0;
      regVec_2548 <= 8'h0;
      regVec_2549 <= 8'h0;
      regVec_2550 <= 8'h0;
      regVec_2551 <= 8'h0;
      regVec_2552 <= 8'h0;
      regVec_2553 <= 8'h0;
      regVec_2554 <= 8'h0;
      regVec_2555 <= 8'h0;
      regVec_2556 <= 8'h0;
      regVec_2557 <= 8'h0;
      regVec_2558 <= 8'h0;
      regVec_2559 <= 8'h0;
      regVec_2560 <= 8'h0;
      regVec_2561 <= 8'h0;
      regVec_2562 <= 8'h0;
      regVec_2563 <= 8'h0;
      regVec_2564 <= 8'h0;
      regVec_2565 <= 8'h0;
      regVec_2566 <= 8'h0;
      regVec_2567 <= 8'h0;
      regVec_2568 <= 8'h0;
      regVec_2569 <= 8'h0;
      regVec_2570 <= 8'h0;
      regVec_2571 <= 8'h0;
      regVec_2572 <= 8'h0;
      regVec_2573 <= 8'h0;
      regVec_2574 <= 8'h0;
      regVec_2575 <= 8'h0;
      regVec_2576 <= 8'h0;
      regVec_2577 <= 8'h0;
      regVec_2578 <= 8'h0;
      regVec_2579 <= 8'h0;
      regVec_2580 <= 8'h0;
      regVec_2581 <= 8'h0;
      regVec_2582 <= 8'h0;
      regVec_2583 <= 8'h0;
      regVec_2584 <= 8'h0;
      regVec_2585 <= 8'h0;
      regVec_2586 <= 8'h0;
      regVec_2587 <= 8'h0;
      regVec_2588 <= 8'h0;
      regVec_2589 <= 8'h0;
      regVec_2590 <= 8'h0;
      regVec_2591 <= 8'h0;
      regVec_2592 <= 8'h0;
      regVec_2593 <= 8'h0;
      regVec_2594 <= 8'h0;
      regVec_2595 <= 8'h0;
      regVec_2596 <= 8'h0;
      regVec_2597 <= 8'h0;
      regVec_2598 <= 8'h0;
      regVec_2599 <= 8'h0;
      regVec_2600 <= 8'h0;
      regVec_2601 <= 8'h0;
      regVec_2602 <= 8'h0;
      regVec_2603 <= 8'h0;
      regVec_2604 <= 8'h0;
      regVec_2605 <= 8'h0;
      regVec_2606 <= 8'h0;
      regVec_2607 <= 8'h0;
      regVec_2608 <= 8'h0;
      regVec_2609 <= 8'h0;
      regVec_2610 <= 8'h0;
      regVec_2611 <= 8'h0;
      regVec_2612 <= 8'h0;
      regVec_2613 <= 8'h0;
      regVec_2614 <= 8'h0;
      regVec_2615 <= 8'h0;
      regVec_2616 <= 8'h0;
      regVec_2617 <= 8'h0;
      regVec_2618 <= 8'h0;
      regVec_2619 <= 8'h0;
      regVec_2620 <= 8'h0;
      regVec_2621 <= 8'h0;
      regVec_2622 <= 8'h0;
      regVec_2623 <= 8'h0;
      regVec_2624 <= 8'h0;
      regVec_2625 <= 8'h0;
      regVec_2626 <= 8'h0;
      regVec_2627 <= 8'h0;
      regVec_2628 <= 8'h0;
      regVec_2629 <= 8'h0;
      regVec_2630 <= 8'h0;
      regVec_2631 <= 8'h0;
      regVec_2632 <= 8'h0;
      regVec_2633 <= 8'h0;
      regVec_2634 <= 8'h0;
      regVec_2635 <= 8'h0;
      regVec_2636 <= 8'h0;
      regVec_2637 <= 8'h0;
      regVec_2638 <= 8'h0;
      regVec_2639 <= 8'h0;
      regVec_2640 <= 8'h0;
      regVec_2641 <= 8'h0;
      regVec_2642 <= 8'h0;
      regVec_2643 <= 8'h0;
      regVec_2644 <= 8'h0;
      regVec_2645 <= 8'h0;
      regVec_2646 <= 8'h0;
      regVec_2647 <= 8'h0;
      regVec_2648 <= 8'h0;
      regVec_2649 <= 8'h0;
      regVec_2650 <= 8'h0;
      regVec_2651 <= 8'h0;
      regVec_2652 <= 8'h0;
      regVec_2653 <= 8'h0;
      regVec_2654 <= 8'h0;
      regVec_2655 <= 8'h0;
      regVec_2656 <= 8'h0;
      regVec_2657 <= 8'h0;
      regVec_2658 <= 8'h0;
      regVec_2659 <= 8'h0;
      regVec_2660 <= 8'h0;
      regVec_2661 <= 8'h0;
      regVec_2662 <= 8'h0;
      regVec_2663 <= 8'h0;
      regVec_2664 <= 8'h0;
      regVec_2665 <= 8'h0;
      regVec_2666 <= 8'h0;
      regVec_2667 <= 8'h0;
      regVec_2668 <= 8'h0;
      regVec_2669 <= 8'h0;
      regVec_2670 <= 8'h0;
      regVec_2671 <= 8'h0;
      regVec_2672 <= 8'h0;
      regVec_2673 <= 8'h0;
      regVec_2674 <= 8'h0;
      regVec_2675 <= 8'h0;
      regVec_2676 <= 8'h0;
      regVec_2677 <= 8'h0;
      regVec_2678 <= 8'h0;
      regVec_2679 <= 8'h0;
      regVec_2680 <= 8'h0;
      regVec_2681 <= 8'h0;
      regVec_2682 <= 8'h0;
      regVec_2683 <= 8'h0;
      regVec_2684 <= 8'h0;
      regVec_2685 <= 8'h0;
      regVec_2686 <= 8'h0;
      regVec_2687 <= 8'h0;
      regVec_2688 <= 8'h0;
      regVec_2689 <= 8'h0;
      regVec_2690 <= 8'h0;
      regVec_2691 <= 8'h0;
      regVec_2692 <= 8'h0;
      regVec_2693 <= 8'h0;
      regVec_2694 <= 8'h0;
      regVec_2695 <= 8'h0;
      regVec_2696 <= 8'h0;
      regVec_2697 <= 8'h0;
      regVec_2698 <= 8'h0;
      regVec_2699 <= 8'h0;
      regVec_2700 <= 8'h0;
      regVec_2701 <= 8'h0;
      regVec_2702 <= 8'h0;
      regVec_2703 <= 8'h0;
      regVec_2704 <= 8'h0;
      regVec_2705 <= 8'h0;
      regVec_2706 <= 8'h0;
      regVec_2707 <= 8'h0;
      regVec_2708 <= 8'h0;
      regVec_2709 <= 8'h0;
      regVec_2710 <= 8'h0;
      regVec_2711 <= 8'h0;
      regVec_2712 <= 8'h0;
      regVec_2713 <= 8'h0;
      regVec_2714 <= 8'h0;
      regVec_2715 <= 8'h0;
      regVec_2716 <= 8'h0;
      regVec_2717 <= 8'h0;
      regVec_2718 <= 8'h0;
      regVec_2719 <= 8'h0;
      regVec_2720 <= 8'h0;
      regVec_2721 <= 8'h0;
      regVec_2722 <= 8'h0;
      regVec_2723 <= 8'h0;
      regVec_2724 <= 8'h0;
      regVec_2725 <= 8'h0;
      regVec_2726 <= 8'h0;
      regVec_2727 <= 8'h0;
      regVec_2728 <= 8'h0;
      regVec_2729 <= 8'h0;
      regVec_2730 <= 8'h0;
      regVec_2731 <= 8'h0;
      regVec_2732 <= 8'h0;
      regVec_2733 <= 8'h0;
      regVec_2734 <= 8'h0;
      regVec_2735 <= 8'h0;
      regVec_2736 <= 8'h0;
      regVec_2737 <= 8'h0;
      regVec_2738 <= 8'h0;
      regVec_2739 <= 8'h0;
      regVec_2740 <= 8'h0;
      regVec_2741 <= 8'h0;
      regVec_2742 <= 8'h0;
      regVec_2743 <= 8'h0;
      regVec_2744 <= 8'h0;
      regVec_2745 <= 8'h0;
      regVec_2746 <= 8'h0;
      regVec_2747 <= 8'h0;
      regVec_2748 <= 8'h0;
      regVec_2749 <= 8'h0;
      regVec_2750 <= 8'h0;
      regVec_2751 <= 8'h0;
      regVec_2752 <= 8'h0;
      regVec_2753 <= 8'h0;
      regVec_2754 <= 8'h0;
      regVec_2755 <= 8'h0;
      regVec_2756 <= 8'h0;
      regVec_2757 <= 8'h0;
      regVec_2758 <= 8'h0;
      regVec_2759 <= 8'h0;
      regVec_2760 <= 8'h0;
      regVec_2761 <= 8'h0;
      regVec_2762 <= 8'h0;
      regVec_2763 <= 8'h0;
      regVec_2764 <= 8'h0;
      regVec_2765 <= 8'h0;
      regVec_2766 <= 8'h0;
      regVec_2767 <= 8'h0;
      regVec_2768 <= 8'h0;
      regVec_2769 <= 8'h0;
      regVec_2770 <= 8'h0;
      regVec_2771 <= 8'h0;
      regVec_2772 <= 8'h0;
      regVec_2773 <= 8'h0;
      regVec_2774 <= 8'h0;
      regVec_2775 <= 8'h0;
      regVec_2776 <= 8'h0;
      regVec_2777 <= 8'h0;
      regVec_2778 <= 8'h0;
      regVec_2779 <= 8'h0;
      regVec_2780 <= 8'h0;
      regVec_2781 <= 8'h0;
      regVec_2782 <= 8'h0;
      regVec_2783 <= 8'h0;
      regVec_2784 <= 8'h0;
      regVec_2785 <= 8'h0;
      regVec_2786 <= 8'h0;
      regVec_2787 <= 8'h0;
      regVec_2788 <= 8'h0;
      regVec_2789 <= 8'h0;
      regVec_2790 <= 8'h0;
      regVec_2791 <= 8'h0;
      regVec_2792 <= 8'h0;
      regVec_2793 <= 8'h0;
      regVec_2794 <= 8'h0;
      regVec_2795 <= 8'h0;
      regVec_2796 <= 8'h0;
      regVec_2797 <= 8'h0;
      regVec_2798 <= 8'h0;
      regVec_2799 <= 8'h0;
      regVec_2800 <= 8'h0;
      regVec_2801 <= 8'h0;
      regVec_2802 <= 8'h0;
      regVec_2803 <= 8'h0;
      regVec_2804 <= 8'h0;
      regVec_2805 <= 8'h0;
      regVec_2806 <= 8'h0;
      regVec_2807 <= 8'h0;
      regVec_2808 <= 8'h0;
      regVec_2809 <= 8'h0;
      regVec_2810 <= 8'h0;
      regVec_2811 <= 8'h0;
      regVec_2812 <= 8'h0;
      regVec_2813 <= 8'h0;
      regVec_2814 <= 8'h0;
      regVec_2815 <= 8'h0;
      regVec_2816 <= 8'h0;
      regVec_2817 <= 8'h0;
      regVec_2818 <= 8'h0;
      regVec_2819 <= 8'h0;
      regVec_2820 <= 8'h0;
      regVec_2821 <= 8'h0;
      regVec_2822 <= 8'h0;
      regVec_2823 <= 8'h0;
      regVec_2824 <= 8'h0;
      regVec_2825 <= 8'h0;
      regVec_2826 <= 8'h0;
      regVec_2827 <= 8'h0;
      regVec_2828 <= 8'h0;
      regVec_2829 <= 8'h0;
      regVec_2830 <= 8'h0;
      regVec_2831 <= 8'h0;
      regVec_2832 <= 8'h0;
      regVec_2833 <= 8'h0;
      regVec_2834 <= 8'h0;
      regVec_2835 <= 8'h0;
      regVec_2836 <= 8'h0;
      regVec_2837 <= 8'h0;
      regVec_2838 <= 8'h0;
      regVec_2839 <= 8'h0;
      regVec_2840 <= 8'h0;
      regVec_2841 <= 8'h0;
      regVec_2842 <= 8'h0;
      regVec_2843 <= 8'h0;
      regVec_2844 <= 8'h0;
      regVec_2845 <= 8'h0;
      regVec_2846 <= 8'h0;
      regVec_2847 <= 8'h0;
      regVec_2848 <= 8'h0;
      regVec_2849 <= 8'h0;
      regVec_2850 <= 8'h0;
      regVec_2851 <= 8'h0;
      regVec_2852 <= 8'h0;
      regVec_2853 <= 8'h0;
      regVec_2854 <= 8'h0;
      regVec_2855 <= 8'h0;
      regVec_2856 <= 8'h0;
      regVec_2857 <= 8'h0;
      regVec_2858 <= 8'h0;
      regVec_2859 <= 8'h0;
      regVec_2860 <= 8'h0;
      regVec_2861 <= 8'h0;
      regVec_2862 <= 8'h0;
      regVec_2863 <= 8'h0;
      regVec_2864 <= 8'h0;
      regVec_2865 <= 8'h0;
      regVec_2866 <= 8'h0;
      regVec_2867 <= 8'h0;
      regVec_2868 <= 8'h0;
      regVec_2869 <= 8'h0;
      regVec_2870 <= 8'h0;
      regVec_2871 <= 8'h0;
      regVec_2872 <= 8'h0;
      regVec_2873 <= 8'h0;
      regVec_2874 <= 8'h0;
      regVec_2875 <= 8'h0;
      regVec_2876 <= 8'h0;
      regVec_2877 <= 8'h0;
      regVec_2878 <= 8'h0;
      regVec_2879 <= 8'h0;
      regVec_2880 <= 8'h0;
      regVec_2881 <= 8'h0;
      regVec_2882 <= 8'h0;
      regVec_2883 <= 8'h0;
      regVec_2884 <= 8'h0;
      regVec_2885 <= 8'h0;
      regVec_2886 <= 8'h0;
      regVec_2887 <= 8'h0;
      regVec_2888 <= 8'h0;
      regVec_2889 <= 8'h0;
      regVec_2890 <= 8'h0;
      regVec_2891 <= 8'h0;
      regVec_2892 <= 8'h0;
      regVec_2893 <= 8'h0;
      regVec_2894 <= 8'h0;
      regVec_2895 <= 8'h0;
      regVec_2896 <= 8'h0;
      regVec_2897 <= 8'h0;
      regVec_2898 <= 8'h0;
      regVec_2899 <= 8'h0;
      regVec_2900 <= 8'h0;
      regVec_2901 <= 8'h0;
      regVec_2902 <= 8'h0;
      regVec_2903 <= 8'h0;
      regVec_2904 <= 8'h0;
      regVec_2905 <= 8'h0;
      regVec_2906 <= 8'h0;
      regVec_2907 <= 8'h0;
      regVec_2908 <= 8'h0;
      regVec_2909 <= 8'h0;
      regVec_2910 <= 8'h0;
      regVec_2911 <= 8'h0;
      regVec_2912 <= 8'h0;
      regVec_2913 <= 8'h0;
      regVec_2914 <= 8'h0;
      regVec_2915 <= 8'h0;
      regVec_2916 <= 8'h0;
      regVec_2917 <= 8'h0;
      regVec_2918 <= 8'h0;
      regVec_2919 <= 8'h0;
      regVec_2920 <= 8'h0;
      regVec_2921 <= 8'h0;
      regVec_2922 <= 8'h0;
      regVec_2923 <= 8'h0;
      regVec_2924 <= 8'h0;
      regVec_2925 <= 8'h0;
      regVec_2926 <= 8'h0;
      regVec_2927 <= 8'h0;
      regVec_2928 <= 8'h0;
      regVec_2929 <= 8'h0;
      regVec_2930 <= 8'h0;
      regVec_2931 <= 8'h0;
      regVec_2932 <= 8'h0;
      regVec_2933 <= 8'h0;
      regVec_2934 <= 8'h0;
      regVec_2935 <= 8'h0;
      regVec_2936 <= 8'h0;
      regVec_2937 <= 8'h0;
      regVec_2938 <= 8'h0;
      regVec_2939 <= 8'h0;
      regVec_2940 <= 8'h0;
      regVec_2941 <= 8'h0;
      regVec_2942 <= 8'h0;
      regVec_2943 <= 8'h0;
      regVec_2944 <= 8'h0;
      regVec_2945 <= 8'h0;
      regVec_2946 <= 8'h0;
      regVec_2947 <= 8'h0;
      regVec_2948 <= 8'h0;
      regVec_2949 <= 8'h0;
      regVec_2950 <= 8'h0;
      regVec_2951 <= 8'h0;
      regVec_2952 <= 8'h0;
      regVec_2953 <= 8'h0;
      regVec_2954 <= 8'h0;
      regVec_2955 <= 8'h0;
      regVec_2956 <= 8'h0;
      regVec_2957 <= 8'h0;
      regVec_2958 <= 8'h0;
      regVec_2959 <= 8'h0;
      regVec_2960 <= 8'h0;
      regVec_2961 <= 8'h0;
      regVec_2962 <= 8'h0;
      regVec_2963 <= 8'h0;
      regVec_2964 <= 8'h0;
      regVec_2965 <= 8'h0;
      regVec_2966 <= 8'h0;
      regVec_2967 <= 8'h0;
      regVec_2968 <= 8'h0;
      regVec_2969 <= 8'h0;
      regVec_2970 <= 8'h0;
      regVec_2971 <= 8'h0;
      regVec_2972 <= 8'h0;
      regVec_2973 <= 8'h0;
      regVec_2974 <= 8'h0;
      regVec_2975 <= 8'h0;
      regVec_2976 <= 8'h0;
      regVec_2977 <= 8'h0;
      regVec_2978 <= 8'h0;
      regVec_2979 <= 8'h0;
      regVec_2980 <= 8'h0;
      regVec_2981 <= 8'h0;
      regVec_2982 <= 8'h0;
      regVec_2983 <= 8'h0;
      regVec_2984 <= 8'h0;
      regVec_2985 <= 8'h0;
      regVec_2986 <= 8'h0;
      regVec_2987 <= 8'h0;
      regVec_2988 <= 8'h0;
      regVec_2989 <= 8'h0;
      regVec_2990 <= 8'h0;
      regVec_2991 <= 8'h0;
      regVec_2992 <= 8'h0;
      regVec_2993 <= 8'h0;
      regVec_2994 <= 8'h0;
      regVec_2995 <= 8'h0;
      regVec_2996 <= 8'h0;
      regVec_2997 <= 8'h0;
      regVec_2998 <= 8'h0;
      regVec_2999 <= 8'h0;
      regVec_3000 <= 8'h0;
      regVec_3001 <= 8'h0;
      regVec_3002 <= 8'h0;
      regVec_3003 <= 8'h0;
      regVec_3004 <= 8'h0;
      regVec_3005 <= 8'h0;
      regVec_3006 <= 8'h0;
      regVec_3007 <= 8'h0;
      regVec_3008 <= 8'h0;
      regVec_3009 <= 8'h0;
      regVec_3010 <= 8'h0;
      regVec_3011 <= 8'h0;
      regVec_3012 <= 8'h0;
      regVec_3013 <= 8'h0;
      regVec_3014 <= 8'h0;
      regVec_3015 <= 8'h0;
      regVec_3016 <= 8'h0;
      regVec_3017 <= 8'h0;
      regVec_3018 <= 8'h0;
      regVec_3019 <= 8'h0;
      regVec_3020 <= 8'h0;
      regVec_3021 <= 8'h0;
      regVec_3022 <= 8'h0;
      regVec_3023 <= 8'h0;
      regVec_3024 <= 8'h0;
      regVec_3025 <= 8'h0;
      regVec_3026 <= 8'h0;
      regVec_3027 <= 8'h0;
      regVec_3028 <= 8'h0;
      regVec_3029 <= 8'h0;
      regVec_3030 <= 8'h0;
      regVec_3031 <= 8'h0;
      regVec_3032 <= 8'h0;
      regVec_3033 <= 8'h0;
      regVec_3034 <= 8'h0;
      regVec_3035 <= 8'h0;
      regVec_3036 <= 8'h0;
      regVec_3037 <= 8'h0;
      regVec_3038 <= 8'h0;
      regVec_3039 <= 8'h0;
      regVec_3040 <= 8'h0;
      regVec_3041 <= 8'h0;
      regVec_3042 <= 8'h0;
      regVec_3043 <= 8'h0;
      regVec_3044 <= 8'h0;
      regVec_3045 <= 8'h0;
      regVec_3046 <= 8'h0;
      regVec_3047 <= 8'h0;
      regVec_3048 <= 8'h0;
      regVec_3049 <= 8'h0;
      regVec_3050 <= 8'h0;
      regVec_3051 <= 8'h0;
      regVec_3052 <= 8'h0;
      regVec_3053 <= 8'h0;
      regVec_3054 <= 8'h0;
      regVec_3055 <= 8'h0;
      regVec_3056 <= 8'h0;
      regVec_3057 <= 8'h0;
      regVec_3058 <= 8'h0;
      regVec_3059 <= 8'h0;
      regVec_3060 <= 8'h0;
      regVec_3061 <= 8'h0;
      regVec_3062 <= 8'h0;
      regVec_3063 <= 8'h0;
      regVec_3064 <= 8'h0;
      regVec_3065 <= 8'h0;
      regVec_3066 <= 8'h0;
      regVec_3067 <= 8'h0;
      regVec_3068 <= 8'h0;
      regVec_3069 <= 8'h0;
      regVec_3070 <= 8'h0;
      regVec_3071 <= 8'h0;
      regVec_3072 <= 8'h0;
      regVec_3073 <= 8'h0;
      regVec_3074 <= 8'h0;
      regVec_3075 <= 8'h0;
      regVec_3076 <= 8'h0;
      regVec_3077 <= 8'h0;
      regVec_3078 <= 8'h0;
      regVec_3079 <= 8'h0;
      regVec_3080 <= 8'h0;
      regVec_3081 <= 8'h0;
      regVec_3082 <= 8'h0;
      regVec_3083 <= 8'h0;
      regVec_3084 <= 8'h0;
      regVec_3085 <= 8'h0;
      regVec_3086 <= 8'h0;
      regVec_3087 <= 8'h0;
      regVec_3088 <= 8'h0;
      regVec_3089 <= 8'h0;
      regVec_3090 <= 8'h0;
      regVec_3091 <= 8'h0;
      regVec_3092 <= 8'h0;
      regVec_3093 <= 8'h0;
      regVec_3094 <= 8'h0;
      regVec_3095 <= 8'h0;
      regVec_3096 <= 8'h0;
      regVec_3097 <= 8'h0;
      regVec_3098 <= 8'h0;
      regVec_3099 <= 8'h0;
      regVec_3100 <= 8'h0;
      regVec_3101 <= 8'h0;
      regVec_3102 <= 8'h0;
      regVec_3103 <= 8'h0;
      regVec_3104 <= 8'h0;
      regVec_3105 <= 8'h0;
      regVec_3106 <= 8'h0;
      regVec_3107 <= 8'h0;
      regVec_3108 <= 8'h0;
      regVec_3109 <= 8'h0;
      regVec_3110 <= 8'h0;
      regVec_3111 <= 8'h0;
      regVec_3112 <= 8'h0;
      regVec_3113 <= 8'h0;
      regVec_3114 <= 8'h0;
      regVec_3115 <= 8'h0;
      regVec_3116 <= 8'h0;
      regVec_3117 <= 8'h0;
      regVec_3118 <= 8'h0;
      regVec_3119 <= 8'h0;
      regVec_3120 <= 8'h0;
      regVec_3121 <= 8'h0;
      regVec_3122 <= 8'h0;
      regVec_3123 <= 8'h0;
      regVec_3124 <= 8'h0;
      regVec_3125 <= 8'h0;
      regVec_3126 <= 8'h0;
      regVec_3127 <= 8'h0;
      regVec_3128 <= 8'h0;
      regVec_3129 <= 8'h0;
      regVec_3130 <= 8'h0;
      regVec_3131 <= 8'h0;
      regVec_3132 <= 8'h0;
      regVec_3133 <= 8'h0;
      regVec_3134 <= 8'h0;
      regVec_3135 <= 8'h0;
      regVec_3136 <= 8'h0;
      regVec_3137 <= 8'h0;
      regVec_3138 <= 8'h0;
      regVec_3139 <= 8'h0;
      regVec_3140 <= 8'h0;
      regVec_3141 <= 8'h0;
      regVec_3142 <= 8'h0;
      regVec_3143 <= 8'h0;
      regVec_3144 <= 8'h0;
      regVec_3145 <= 8'h0;
      regVec_3146 <= 8'h0;
      regVec_3147 <= 8'h0;
      regVec_3148 <= 8'h0;
      regVec_3149 <= 8'h0;
      regVec_3150 <= 8'h0;
      regVec_3151 <= 8'h0;
      regVec_3152 <= 8'h0;
      regVec_3153 <= 8'h0;
      regVec_3154 <= 8'h0;
      regVec_3155 <= 8'h0;
      regVec_3156 <= 8'h0;
      regVec_3157 <= 8'h0;
      regVec_3158 <= 8'h0;
      regVec_3159 <= 8'h0;
      regVec_3160 <= 8'h0;
      regVec_3161 <= 8'h0;
      regVec_3162 <= 8'h0;
      regVec_3163 <= 8'h0;
      regVec_3164 <= 8'h0;
      regVec_3165 <= 8'h0;
      regVec_3166 <= 8'h0;
      regVec_3167 <= 8'h0;
      regVec_3168 <= 8'h0;
      regVec_3169 <= 8'h0;
      regVec_3170 <= 8'h0;
      regVec_3171 <= 8'h0;
      regVec_3172 <= 8'h0;
      regVec_3173 <= 8'h0;
      regVec_3174 <= 8'h0;
      regVec_3175 <= 8'h0;
      regVec_3176 <= 8'h0;
      regVec_3177 <= 8'h0;
      regVec_3178 <= 8'h0;
      regVec_3179 <= 8'h0;
      regVec_3180 <= 8'h0;
      regVec_3181 <= 8'h0;
      regVec_3182 <= 8'h0;
      regVec_3183 <= 8'h0;
      regVec_3184 <= 8'h0;
      regVec_3185 <= 8'h0;
      regVec_3186 <= 8'h0;
      regVec_3187 <= 8'h0;
      regVec_3188 <= 8'h0;
      regVec_3189 <= 8'h0;
      regVec_3190 <= 8'h0;
      regVec_3191 <= 8'h0;
      regVec_3192 <= 8'h0;
      regVec_3193 <= 8'h0;
      regVec_3194 <= 8'h0;
      regVec_3195 <= 8'h0;
      regVec_3196 <= 8'h0;
      regVec_3197 <= 8'h0;
      regVec_3198 <= 8'h0;
      regVec_3199 <= 8'h0;
      regVec_3200 <= 8'h0;
      regVec_3201 <= 8'h0;
      regVec_3202 <= 8'h0;
      regVec_3203 <= 8'h0;
      regVec_3204 <= 8'h0;
      regVec_3205 <= 8'h0;
      regVec_3206 <= 8'h0;
      regVec_3207 <= 8'h0;
      regVec_3208 <= 8'h0;
      regVec_3209 <= 8'h0;
      regVec_3210 <= 8'h0;
      regVec_3211 <= 8'h0;
      regVec_3212 <= 8'h0;
      regVec_3213 <= 8'h0;
      regVec_3214 <= 8'h0;
      regVec_3215 <= 8'h0;
      regVec_3216 <= 8'h0;
      regVec_3217 <= 8'h0;
      regVec_3218 <= 8'h0;
      regVec_3219 <= 8'h0;
      regVec_3220 <= 8'h0;
      regVec_3221 <= 8'h0;
      regVec_3222 <= 8'h0;
      regVec_3223 <= 8'h0;
      regVec_3224 <= 8'h0;
      regVec_3225 <= 8'h0;
      regVec_3226 <= 8'h0;
      regVec_3227 <= 8'h0;
      regVec_3228 <= 8'h0;
      regVec_3229 <= 8'h0;
      regVec_3230 <= 8'h0;
      regVec_3231 <= 8'h0;
      regVec_3232 <= 8'h0;
      regVec_3233 <= 8'h0;
      regVec_3234 <= 8'h0;
      regVec_3235 <= 8'h0;
      regVec_3236 <= 8'h0;
      regVec_3237 <= 8'h0;
      regVec_3238 <= 8'h0;
      regVec_3239 <= 8'h0;
      regVec_3240 <= 8'h0;
      regVec_3241 <= 8'h0;
      regVec_3242 <= 8'h0;
      regVec_3243 <= 8'h0;
      regVec_3244 <= 8'h0;
      regVec_3245 <= 8'h0;
      regVec_3246 <= 8'h0;
      regVec_3247 <= 8'h0;
      regVec_3248 <= 8'h0;
      regVec_3249 <= 8'h0;
      regVec_3250 <= 8'h0;
      regVec_3251 <= 8'h0;
      regVec_3252 <= 8'h0;
      regVec_3253 <= 8'h0;
      regVec_3254 <= 8'h0;
      regVec_3255 <= 8'h0;
      regVec_3256 <= 8'h0;
      regVec_3257 <= 8'h0;
      regVec_3258 <= 8'h0;
      regVec_3259 <= 8'h0;
      regVec_3260 <= 8'h0;
      regVec_3261 <= 8'h0;
      regVec_3262 <= 8'h0;
      regVec_3263 <= 8'h0;
      regVec_3264 <= 8'h0;
      regVec_3265 <= 8'h0;
      regVec_3266 <= 8'h0;
      regVec_3267 <= 8'h0;
      regVec_3268 <= 8'h0;
      regVec_3269 <= 8'h0;
      regVec_3270 <= 8'h0;
      regVec_3271 <= 8'h0;
      regVec_3272 <= 8'h0;
      regVec_3273 <= 8'h0;
      regVec_3274 <= 8'h0;
      regVec_3275 <= 8'h0;
      regVec_3276 <= 8'h0;
      regVec_3277 <= 8'h0;
      regVec_3278 <= 8'h0;
      regVec_3279 <= 8'h0;
      regVec_3280 <= 8'h0;
      regVec_3281 <= 8'h0;
      regVec_3282 <= 8'h0;
      regVec_3283 <= 8'h0;
      regVec_3284 <= 8'h0;
      regVec_3285 <= 8'h0;
      regVec_3286 <= 8'h0;
      regVec_3287 <= 8'h0;
      regVec_3288 <= 8'h0;
      regVec_3289 <= 8'h0;
      regVec_3290 <= 8'h0;
      regVec_3291 <= 8'h0;
      regVec_3292 <= 8'h0;
      regVec_3293 <= 8'h0;
      regVec_3294 <= 8'h0;
      regVec_3295 <= 8'h0;
      regVec_3296 <= 8'h0;
      regVec_3297 <= 8'h0;
      regVec_3298 <= 8'h0;
      regVec_3299 <= 8'h0;
      regVec_3300 <= 8'h0;
      regVec_3301 <= 8'h0;
      regVec_3302 <= 8'h0;
      regVec_3303 <= 8'h0;
      regVec_3304 <= 8'h0;
      regVec_3305 <= 8'h0;
      regVec_3306 <= 8'h0;
      regVec_3307 <= 8'h0;
      regVec_3308 <= 8'h0;
      regVec_3309 <= 8'h0;
      regVec_3310 <= 8'h0;
      regVec_3311 <= 8'h0;
      regVec_3312 <= 8'h0;
      regVec_3313 <= 8'h0;
      regVec_3314 <= 8'h0;
      regVec_3315 <= 8'h0;
      regVec_3316 <= 8'h0;
      regVec_3317 <= 8'h0;
      regVec_3318 <= 8'h0;
      regVec_3319 <= 8'h0;
      regVec_3320 <= 8'h0;
      regVec_3321 <= 8'h0;
      regVec_3322 <= 8'h0;
      regVec_3323 <= 8'h0;
      regVec_3324 <= 8'h0;
      regVec_3325 <= 8'h0;
      regVec_3326 <= 8'h0;
      regVec_3327 <= 8'h0;
      regVec_3328 <= 8'h0;
      regVec_3329 <= 8'h0;
      regVec_3330 <= 8'h0;
      regVec_3331 <= 8'h0;
      regVec_3332 <= 8'h0;
      regVec_3333 <= 8'h0;
      regVec_3334 <= 8'h0;
      regVec_3335 <= 8'h0;
      regVec_3336 <= 8'h0;
      regVec_3337 <= 8'h0;
      regVec_3338 <= 8'h0;
      regVec_3339 <= 8'h0;
      regVec_3340 <= 8'h0;
      regVec_3341 <= 8'h0;
      regVec_3342 <= 8'h0;
      regVec_3343 <= 8'h0;
      regVec_3344 <= 8'h0;
      regVec_3345 <= 8'h0;
      regVec_3346 <= 8'h0;
      regVec_3347 <= 8'h0;
      regVec_3348 <= 8'h0;
      regVec_3349 <= 8'h0;
      regVec_3350 <= 8'h0;
      regVec_3351 <= 8'h0;
      regVec_3352 <= 8'h0;
      regVec_3353 <= 8'h0;
      regVec_3354 <= 8'h0;
      regVec_3355 <= 8'h0;
      regVec_3356 <= 8'h0;
      regVec_3357 <= 8'h0;
      regVec_3358 <= 8'h0;
      regVec_3359 <= 8'h0;
      regVec_3360 <= 8'h0;
      regVec_3361 <= 8'h0;
      regVec_3362 <= 8'h0;
      regVec_3363 <= 8'h0;
      regVec_3364 <= 8'h0;
      regVec_3365 <= 8'h0;
      regVec_3366 <= 8'h0;
      regVec_3367 <= 8'h0;
      regVec_3368 <= 8'h0;
      regVec_3369 <= 8'h0;
      regVec_3370 <= 8'h0;
      regVec_3371 <= 8'h0;
      regVec_3372 <= 8'h0;
      regVec_3373 <= 8'h0;
      regVec_3374 <= 8'h0;
      regVec_3375 <= 8'h0;
      regVec_3376 <= 8'h0;
      regVec_3377 <= 8'h0;
      regVec_3378 <= 8'h0;
      regVec_3379 <= 8'h0;
      regVec_3380 <= 8'h0;
      regVec_3381 <= 8'h0;
      regVec_3382 <= 8'h0;
      regVec_3383 <= 8'h0;
      regVec_3384 <= 8'h0;
      regVec_3385 <= 8'h0;
      regVec_3386 <= 8'h0;
      regVec_3387 <= 8'h0;
      regVec_3388 <= 8'h0;
      regVec_3389 <= 8'h0;
      regVec_3390 <= 8'h0;
      regVec_3391 <= 8'h0;
      regVec_3392 <= 8'h0;
      regVec_3393 <= 8'h0;
      regVec_3394 <= 8'h0;
      regVec_3395 <= 8'h0;
      regVec_3396 <= 8'h0;
      regVec_3397 <= 8'h0;
      regVec_3398 <= 8'h0;
      regVec_3399 <= 8'h0;
      regVec_3400 <= 8'h0;
      regVec_3401 <= 8'h0;
      regVec_3402 <= 8'h0;
      regVec_3403 <= 8'h0;
      regVec_3404 <= 8'h0;
      regVec_3405 <= 8'h0;
      regVec_3406 <= 8'h0;
      regVec_3407 <= 8'h0;
      regVec_3408 <= 8'h0;
      regVec_3409 <= 8'h0;
      regVec_3410 <= 8'h0;
      regVec_3411 <= 8'h0;
      regVec_3412 <= 8'h0;
      regVec_3413 <= 8'h0;
      regVec_3414 <= 8'h0;
      regVec_3415 <= 8'h0;
      regVec_3416 <= 8'h0;
      regVec_3417 <= 8'h0;
      regVec_3418 <= 8'h0;
      regVec_3419 <= 8'h0;
      regVec_3420 <= 8'h0;
      regVec_3421 <= 8'h0;
      regVec_3422 <= 8'h0;
      regVec_3423 <= 8'h0;
      regVec_3424 <= 8'h0;
      regVec_3425 <= 8'h0;
      regVec_3426 <= 8'h0;
      regVec_3427 <= 8'h0;
      regVec_3428 <= 8'h0;
      regVec_3429 <= 8'h0;
      regVec_3430 <= 8'h0;
      regVec_3431 <= 8'h0;
      regVec_3432 <= 8'h0;
      regVec_3433 <= 8'h0;
      regVec_3434 <= 8'h0;
      regVec_3435 <= 8'h0;
      regVec_3436 <= 8'h0;
      regVec_3437 <= 8'h0;
      regVec_3438 <= 8'h0;
      regVec_3439 <= 8'h0;
      regVec_3440 <= 8'h0;
      regVec_3441 <= 8'h0;
      regVec_3442 <= 8'h0;
      regVec_3443 <= 8'h0;
      regVec_3444 <= 8'h0;
      regVec_3445 <= 8'h0;
      regVec_3446 <= 8'h0;
      regVec_3447 <= 8'h0;
      regVec_3448 <= 8'h0;
      regVec_3449 <= 8'h0;
      regVec_3450 <= 8'h0;
      regVec_3451 <= 8'h0;
      regVec_3452 <= 8'h0;
      regVec_3453 <= 8'h0;
      regVec_3454 <= 8'h0;
      regVec_3455 <= 8'h0;
      regVec_3456 <= 8'h0;
      regVec_3457 <= 8'h0;
      regVec_3458 <= 8'h0;
      regVec_3459 <= 8'h0;
      regVec_3460 <= 8'h0;
      regVec_3461 <= 8'h0;
      regVec_3462 <= 8'h0;
      regVec_3463 <= 8'h0;
      regVec_3464 <= 8'h0;
      regVec_3465 <= 8'h0;
      regVec_3466 <= 8'h0;
      regVec_3467 <= 8'h0;
      regVec_3468 <= 8'h0;
      regVec_3469 <= 8'h0;
      regVec_3470 <= 8'h0;
      regVec_3471 <= 8'h0;
      regVec_3472 <= 8'h0;
      regVec_3473 <= 8'h0;
      regVec_3474 <= 8'h0;
      regVec_3475 <= 8'h0;
      regVec_3476 <= 8'h0;
      regVec_3477 <= 8'h0;
      regVec_3478 <= 8'h0;
      regVec_3479 <= 8'h0;
      regVec_3480 <= 8'h0;
      regVec_3481 <= 8'h0;
      regVec_3482 <= 8'h0;
      regVec_3483 <= 8'h0;
      regVec_3484 <= 8'h0;
      regVec_3485 <= 8'h0;
      regVec_3486 <= 8'h0;
      regVec_3487 <= 8'h0;
      regVec_3488 <= 8'h0;
      regVec_3489 <= 8'h0;
      regVec_3490 <= 8'h0;
      regVec_3491 <= 8'h0;
      regVec_3492 <= 8'h0;
      regVec_3493 <= 8'h0;
      regVec_3494 <= 8'h0;
      regVec_3495 <= 8'h0;
      regVec_3496 <= 8'h0;
      regVec_3497 <= 8'h0;
      regVec_3498 <= 8'h0;
      regVec_3499 <= 8'h0;
      regVec_3500 <= 8'h0;
      regVec_3501 <= 8'h0;
      regVec_3502 <= 8'h0;
      regVec_3503 <= 8'h0;
      regVec_3504 <= 8'h0;
      regVec_3505 <= 8'h0;
      regVec_3506 <= 8'h0;
      regVec_3507 <= 8'h0;
      regVec_3508 <= 8'h0;
      regVec_3509 <= 8'h0;
      regVec_3510 <= 8'h0;
      regVec_3511 <= 8'h0;
      regVec_3512 <= 8'h0;
      regVec_3513 <= 8'h0;
      regVec_3514 <= 8'h0;
      regVec_3515 <= 8'h0;
      regVec_3516 <= 8'h0;
      regVec_3517 <= 8'h0;
      regVec_3518 <= 8'h0;
      regVec_3519 <= 8'h0;
      regVec_3520 <= 8'h0;
      regVec_3521 <= 8'h0;
      regVec_3522 <= 8'h0;
      regVec_3523 <= 8'h0;
      regVec_3524 <= 8'h0;
      regVec_3525 <= 8'h0;
      regVec_3526 <= 8'h0;
      regVec_3527 <= 8'h0;
      regVec_3528 <= 8'h0;
      regVec_3529 <= 8'h0;
      regVec_3530 <= 8'h0;
      regVec_3531 <= 8'h0;
      regVec_3532 <= 8'h0;
      regVec_3533 <= 8'h0;
      regVec_3534 <= 8'h0;
      regVec_3535 <= 8'h0;
      regVec_3536 <= 8'h0;
      regVec_3537 <= 8'h0;
      regVec_3538 <= 8'h0;
      regVec_3539 <= 8'h0;
      regVec_3540 <= 8'h0;
      regVec_3541 <= 8'h0;
      regVec_3542 <= 8'h0;
      regVec_3543 <= 8'h0;
      regVec_3544 <= 8'h0;
      regVec_3545 <= 8'h0;
      regVec_3546 <= 8'h0;
      regVec_3547 <= 8'h0;
      regVec_3548 <= 8'h0;
      regVec_3549 <= 8'h0;
      regVec_3550 <= 8'h0;
      regVec_3551 <= 8'h0;
      regVec_3552 <= 8'h0;
      regVec_3553 <= 8'h0;
      regVec_3554 <= 8'h0;
      regVec_3555 <= 8'h0;
      regVec_3556 <= 8'h0;
      regVec_3557 <= 8'h0;
      regVec_3558 <= 8'h0;
      regVec_3559 <= 8'h0;
      regVec_3560 <= 8'h0;
      regVec_3561 <= 8'h0;
      regVec_3562 <= 8'h0;
      regVec_3563 <= 8'h0;
      regVec_3564 <= 8'h0;
      regVec_3565 <= 8'h0;
      regVec_3566 <= 8'h0;
      regVec_3567 <= 8'h0;
      regVec_3568 <= 8'h0;
      regVec_3569 <= 8'h0;
      regVec_3570 <= 8'h0;
      regVec_3571 <= 8'h0;
      regVec_3572 <= 8'h0;
      regVec_3573 <= 8'h0;
      regVec_3574 <= 8'h0;
      regVec_3575 <= 8'h0;
      regVec_3576 <= 8'h0;
      regVec_3577 <= 8'h0;
      regVec_3578 <= 8'h0;
      regVec_3579 <= 8'h0;
      regVec_3580 <= 8'h0;
      regVec_3581 <= 8'h0;
      regVec_3582 <= 8'h0;
      regVec_3583 <= 8'h0;
      regVec_3584 <= 8'h0;
      regVec_3585 <= 8'h0;
      regVec_3586 <= 8'h0;
      regVec_3587 <= 8'h0;
      regVec_3588 <= 8'h0;
      regVec_3589 <= 8'h0;
      regVec_3590 <= 8'h0;
      regVec_3591 <= 8'h0;
      regVec_3592 <= 8'h0;
      regVec_3593 <= 8'h0;
      regVec_3594 <= 8'h0;
      regVec_3595 <= 8'h0;
      regVec_3596 <= 8'h0;
      regVec_3597 <= 8'h0;
      regVec_3598 <= 8'h0;
      regVec_3599 <= 8'h0;
      regVec_3600 <= 8'h0;
      regVec_3601 <= 8'h0;
      regVec_3602 <= 8'h0;
      regVec_3603 <= 8'h0;
      regVec_3604 <= 8'h0;
      regVec_3605 <= 8'h0;
      regVec_3606 <= 8'h0;
      regVec_3607 <= 8'h0;
      regVec_3608 <= 8'h0;
      regVec_3609 <= 8'h0;
      regVec_3610 <= 8'h0;
      regVec_3611 <= 8'h0;
      regVec_3612 <= 8'h0;
      regVec_3613 <= 8'h0;
      regVec_3614 <= 8'h0;
      regVec_3615 <= 8'h0;
      regVec_3616 <= 8'h0;
      regVec_3617 <= 8'h0;
      regVec_3618 <= 8'h0;
      regVec_3619 <= 8'h0;
      regVec_3620 <= 8'h0;
      regVec_3621 <= 8'h0;
      regVec_3622 <= 8'h0;
      regVec_3623 <= 8'h0;
      regVec_3624 <= 8'h0;
      regVec_3625 <= 8'h0;
      regVec_3626 <= 8'h0;
      regVec_3627 <= 8'h0;
      regVec_3628 <= 8'h0;
      regVec_3629 <= 8'h0;
      regVec_3630 <= 8'h0;
      regVec_3631 <= 8'h0;
      regVec_3632 <= 8'h0;
      regVec_3633 <= 8'h0;
      regVec_3634 <= 8'h0;
      regVec_3635 <= 8'h0;
      regVec_3636 <= 8'h0;
      regVec_3637 <= 8'h0;
      regVec_3638 <= 8'h0;
      regVec_3639 <= 8'h0;
      regVec_3640 <= 8'h0;
      regVec_3641 <= 8'h0;
      regVec_3642 <= 8'h0;
      regVec_3643 <= 8'h0;
      regVec_3644 <= 8'h0;
      regVec_3645 <= 8'h0;
      regVec_3646 <= 8'h0;
      regVec_3647 <= 8'h0;
      regVec_3648 <= 8'h0;
      regVec_3649 <= 8'h0;
      regVec_3650 <= 8'h0;
      regVec_3651 <= 8'h0;
      regVec_3652 <= 8'h0;
      regVec_3653 <= 8'h0;
      regVec_3654 <= 8'h0;
      regVec_3655 <= 8'h0;
      regVec_3656 <= 8'h0;
      regVec_3657 <= 8'h0;
      regVec_3658 <= 8'h0;
      regVec_3659 <= 8'h0;
      regVec_3660 <= 8'h0;
      regVec_3661 <= 8'h0;
      regVec_3662 <= 8'h0;
      regVec_3663 <= 8'h0;
      regVec_3664 <= 8'h0;
      regVec_3665 <= 8'h0;
      regVec_3666 <= 8'h0;
      regVec_3667 <= 8'h0;
      regVec_3668 <= 8'h0;
      regVec_3669 <= 8'h0;
      regVec_3670 <= 8'h0;
      regVec_3671 <= 8'h0;
      regVec_3672 <= 8'h0;
      regVec_3673 <= 8'h0;
      regVec_3674 <= 8'h0;
      regVec_3675 <= 8'h0;
      regVec_3676 <= 8'h0;
      regVec_3677 <= 8'h0;
      regVec_3678 <= 8'h0;
      regVec_3679 <= 8'h0;
      regVec_3680 <= 8'h0;
      regVec_3681 <= 8'h0;
      regVec_3682 <= 8'h0;
      regVec_3683 <= 8'h0;
      regVec_3684 <= 8'h0;
      regVec_3685 <= 8'h0;
      regVec_3686 <= 8'h0;
      regVec_3687 <= 8'h0;
      regVec_3688 <= 8'h0;
      regVec_3689 <= 8'h0;
      regVec_3690 <= 8'h0;
      regVec_3691 <= 8'h0;
      regVec_3692 <= 8'h0;
      regVec_3693 <= 8'h0;
      regVec_3694 <= 8'h0;
      regVec_3695 <= 8'h0;
      regVec_3696 <= 8'h0;
      regVec_3697 <= 8'h0;
      regVec_3698 <= 8'h0;
      regVec_3699 <= 8'h0;
      regVec_3700 <= 8'h0;
      regVec_3701 <= 8'h0;
      regVec_3702 <= 8'h0;
      regVec_3703 <= 8'h0;
      regVec_3704 <= 8'h0;
      regVec_3705 <= 8'h0;
      regVec_3706 <= 8'h0;
      regVec_3707 <= 8'h0;
      regVec_3708 <= 8'h0;
      regVec_3709 <= 8'h0;
      regVec_3710 <= 8'h0;
      regVec_3711 <= 8'h0;
      regVec_3712 <= 8'h0;
      regVec_3713 <= 8'h0;
      regVec_3714 <= 8'h0;
      regVec_3715 <= 8'h0;
      regVec_3716 <= 8'h0;
      regVec_3717 <= 8'h0;
      regVec_3718 <= 8'h0;
      regVec_3719 <= 8'h0;
      regVec_3720 <= 8'h0;
      regVec_3721 <= 8'h0;
      regVec_3722 <= 8'h0;
      regVec_3723 <= 8'h0;
      regVec_3724 <= 8'h0;
      regVec_3725 <= 8'h0;
      regVec_3726 <= 8'h0;
      regVec_3727 <= 8'h0;
      regVec_3728 <= 8'h0;
      regVec_3729 <= 8'h0;
      regVec_3730 <= 8'h0;
      regVec_3731 <= 8'h0;
      regVec_3732 <= 8'h0;
      regVec_3733 <= 8'h0;
      regVec_3734 <= 8'h0;
      regVec_3735 <= 8'h0;
      regVec_3736 <= 8'h0;
      regVec_3737 <= 8'h0;
      regVec_3738 <= 8'h0;
      regVec_3739 <= 8'h0;
      regVec_3740 <= 8'h0;
      regVec_3741 <= 8'h0;
      regVec_3742 <= 8'h0;
      regVec_3743 <= 8'h0;
      regVec_3744 <= 8'h0;
      regVec_3745 <= 8'h0;
      regVec_3746 <= 8'h0;
      regVec_3747 <= 8'h0;
      regVec_3748 <= 8'h0;
      regVec_3749 <= 8'h0;
      regVec_3750 <= 8'h0;
      regVec_3751 <= 8'h0;
      regVec_3752 <= 8'h0;
      regVec_3753 <= 8'h0;
      regVec_3754 <= 8'h0;
      regVec_3755 <= 8'h0;
      regVec_3756 <= 8'h0;
      regVec_3757 <= 8'h0;
      regVec_3758 <= 8'h0;
      regVec_3759 <= 8'h0;
      regVec_3760 <= 8'h0;
      regVec_3761 <= 8'h0;
      regVec_3762 <= 8'h0;
      regVec_3763 <= 8'h0;
      regVec_3764 <= 8'h0;
      regVec_3765 <= 8'h0;
      regVec_3766 <= 8'h0;
      regVec_3767 <= 8'h0;
      regVec_3768 <= 8'h0;
      regVec_3769 <= 8'h0;
      regVec_3770 <= 8'h0;
      regVec_3771 <= 8'h0;
      regVec_3772 <= 8'h0;
      regVec_3773 <= 8'h0;
      regVec_3774 <= 8'h0;
      regVec_3775 <= 8'h0;
      regVec_3776 <= 8'h0;
      regVec_3777 <= 8'h0;
      regVec_3778 <= 8'h0;
      regVec_3779 <= 8'h0;
      regVec_3780 <= 8'h0;
      regVec_3781 <= 8'h0;
      regVec_3782 <= 8'h0;
      regVec_3783 <= 8'h0;
      regVec_3784 <= 8'h0;
      regVec_3785 <= 8'h0;
      regVec_3786 <= 8'h0;
      regVec_3787 <= 8'h0;
      regVec_3788 <= 8'h0;
      regVec_3789 <= 8'h0;
      regVec_3790 <= 8'h0;
      regVec_3791 <= 8'h0;
      regVec_3792 <= 8'h0;
      regVec_3793 <= 8'h0;
      regVec_3794 <= 8'h0;
      regVec_3795 <= 8'h0;
      regVec_3796 <= 8'h0;
      regVec_3797 <= 8'h0;
      regVec_3798 <= 8'h0;
      regVec_3799 <= 8'h0;
      regVec_3800 <= 8'h0;
      regVec_3801 <= 8'h0;
      regVec_3802 <= 8'h0;
      regVec_3803 <= 8'h0;
      regVec_3804 <= 8'h0;
      regVec_3805 <= 8'h0;
      regVec_3806 <= 8'h0;
      regVec_3807 <= 8'h0;
      regVec_3808 <= 8'h0;
      regVec_3809 <= 8'h0;
      regVec_3810 <= 8'h0;
      regVec_3811 <= 8'h0;
      regVec_3812 <= 8'h0;
      regVec_3813 <= 8'h0;
      regVec_3814 <= 8'h0;
      regVec_3815 <= 8'h0;
      regVec_3816 <= 8'h0;
      regVec_3817 <= 8'h0;
      regVec_3818 <= 8'h0;
      regVec_3819 <= 8'h0;
      regVec_3820 <= 8'h0;
      regVec_3821 <= 8'h0;
      regVec_3822 <= 8'h0;
      regVec_3823 <= 8'h0;
      regVec_3824 <= 8'h0;
      regVec_3825 <= 8'h0;
      regVec_3826 <= 8'h0;
      regVec_3827 <= 8'h0;
      regVec_3828 <= 8'h0;
      regVec_3829 <= 8'h0;
      regVec_3830 <= 8'h0;
      regVec_3831 <= 8'h0;
      regVec_3832 <= 8'h0;
      regVec_3833 <= 8'h0;
      regVec_3834 <= 8'h0;
      regVec_3835 <= 8'h0;
      regVec_3836 <= 8'h0;
      regVec_3837 <= 8'h0;
      regVec_3838 <= 8'h0;
      regVec_3839 <= 8'h0;
      regVec_3840 <= 8'h0;
      regVec_3841 <= 8'h0;
      regVec_3842 <= 8'h0;
      regVec_3843 <= 8'h0;
      regVec_3844 <= 8'h0;
      regVec_3845 <= 8'h0;
      regVec_3846 <= 8'h0;
      regVec_3847 <= 8'h0;
      regVec_3848 <= 8'h0;
      regVec_3849 <= 8'h0;
      regVec_3850 <= 8'h0;
      regVec_3851 <= 8'h0;
      regVec_3852 <= 8'h0;
      regVec_3853 <= 8'h0;
      regVec_3854 <= 8'h0;
      regVec_3855 <= 8'h0;
      regVec_3856 <= 8'h0;
      regVec_3857 <= 8'h0;
      regVec_3858 <= 8'h0;
      regVec_3859 <= 8'h0;
      regVec_3860 <= 8'h0;
      regVec_3861 <= 8'h0;
      regVec_3862 <= 8'h0;
      regVec_3863 <= 8'h0;
      regVec_3864 <= 8'h0;
      regVec_3865 <= 8'h0;
      regVec_3866 <= 8'h0;
      regVec_3867 <= 8'h0;
      regVec_3868 <= 8'h0;
      regVec_3869 <= 8'h0;
      regVec_3870 <= 8'h0;
      regVec_3871 <= 8'h0;
      regVec_3872 <= 8'h0;
      regVec_3873 <= 8'h0;
      regVec_3874 <= 8'h0;
      regVec_3875 <= 8'h0;
      regVec_3876 <= 8'h0;
      regVec_3877 <= 8'h0;
      regVec_3878 <= 8'h0;
      regVec_3879 <= 8'h0;
      regVec_3880 <= 8'h0;
      regVec_3881 <= 8'h0;
      regVec_3882 <= 8'h0;
      regVec_3883 <= 8'h0;
      regVec_3884 <= 8'h0;
      regVec_3885 <= 8'h0;
      regVec_3886 <= 8'h0;
      regVec_3887 <= 8'h0;
      regVec_3888 <= 8'h0;
      regVec_3889 <= 8'h0;
      regVec_3890 <= 8'h0;
      regVec_3891 <= 8'h0;
      regVec_3892 <= 8'h0;
      regVec_3893 <= 8'h0;
      regVec_3894 <= 8'h0;
      regVec_3895 <= 8'h0;
      regVec_3896 <= 8'h0;
      regVec_3897 <= 8'h0;
      regVec_3898 <= 8'h0;
      regVec_3899 <= 8'h0;
      regVec_3900 <= 8'h0;
      regVec_3901 <= 8'h0;
      regVec_3902 <= 8'h0;
      regVec_3903 <= 8'h0;
      regVec_3904 <= 8'h0;
      regVec_3905 <= 8'h0;
      regVec_3906 <= 8'h0;
      regVec_3907 <= 8'h0;
      regVec_3908 <= 8'h0;
      regVec_3909 <= 8'h0;
      regVec_3910 <= 8'h0;
      regVec_3911 <= 8'h0;
      regVec_3912 <= 8'h0;
      regVec_3913 <= 8'h0;
      regVec_3914 <= 8'h0;
      regVec_3915 <= 8'h0;
      regVec_3916 <= 8'h0;
      regVec_3917 <= 8'h0;
      regVec_3918 <= 8'h0;
      regVec_3919 <= 8'h0;
      regVec_3920 <= 8'h0;
      regVec_3921 <= 8'h0;
      regVec_3922 <= 8'h0;
      regVec_3923 <= 8'h0;
      regVec_3924 <= 8'h0;
      regVec_3925 <= 8'h0;
      regVec_3926 <= 8'h0;
      regVec_3927 <= 8'h0;
      regVec_3928 <= 8'h0;
      regVec_3929 <= 8'h0;
      regVec_3930 <= 8'h0;
      regVec_3931 <= 8'h0;
      regVec_3932 <= 8'h0;
      regVec_3933 <= 8'h0;
      regVec_3934 <= 8'h0;
      regVec_3935 <= 8'h0;
      regVec_3936 <= 8'h0;
      regVec_3937 <= 8'h0;
      regVec_3938 <= 8'h0;
      regVec_3939 <= 8'h0;
      regVec_3940 <= 8'h0;
      regVec_3941 <= 8'h0;
      regVec_3942 <= 8'h0;
      regVec_3943 <= 8'h0;
      regVec_3944 <= 8'h0;
      regVec_3945 <= 8'h0;
      regVec_3946 <= 8'h0;
      regVec_3947 <= 8'h0;
      regVec_3948 <= 8'h0;
      regVec_3949 <= 8'h0;
      regVec_3950 <= 8'h0;
      regVec_3951 <= 8'h0;
      regVec_3952 <= 8'h0;
      regVec_3953 <= 8'h0;
      regVec_3954 <= 8'h0;
      regVec_3955 <= 8'h0;
      regVec_3956 <= 8'h0;
      regVec_3957 <= 8'h0;
      regVec_3958 <= 8'h0;
      regVec_3959 <= 8'h0;
      regVec_3960 <= 8'h0;
      regVec_3961 <= 8'h0;
      regVec_3962 <= 8'h0;
      regVec_3963 <= 8'h0;
      regVec_3964 <= 8'h0;
      regVec_3965 <= 8'h0;
      regVec_3966 <= 8'h0;
      regVec_3967 <= 8'h0;
      regVec_3968 <= 8'h0;
      regVec_3969 <= 8'h0;
      regVec_3970 <= 8'h0;
      regVec_3971 <= 8'h0;
      regVec_3972 <= 8'h0;
      regVec_3973 <= 8'h0;
      regVec_3974 <= 8'h0;
      regVec_3975 <= 8'h0;
      regVec_3976 <= 8'h0;
      regVec_3977 <= 8'h0;
      regVec_3978 <= 8'h0;
      regVec_3979 <= 8'h0;
      regVec_3980 <= 8'h0;
      regVec_3981 <= 8'h0;
      regVec_3982 <= 8'h0;
      regVec_3983 <= 8'h0;
      regVec_3984 <= 8'h0;
      regVec_3985 <= 8'h0;
      regVec_3986 <= 8'h0;
      regVec_3987 <= 8'h0;
      regVec_3988 <= 8'h0;
      regVec_3989 <= 8'h0;
      regVec_3990 <= 8'h0;
      regVec_3991 <= 8'h0;
      regVec_3992 <= 8'h0;
      regVec_3993 <= 8'h0;
      regVec_3994 <= 8'h0;
      regVec_3995 <= 8'h0;
      regVec_3996 <= 8'h0;
      regVec_3997 <= 8'h0;
      regVec_3998 <= 8'h0;
      regVec_3999 <= 8'h0;
      regVec_4000 <= 8'h0;
      regVec_4001 <= 8'h0;
      regVec_4002 <= 8'h0;
      regVec_4003 <= 8'h0;
      regVec_4004 <= 8'h0;
      regVec_4005 <= 8'h0;
      regVec_4006 <= 8'h0;
      regVec_4007 <= 8'h0;
      regVec_4008 <= 8'h0;
      regVec_4009 <= 8'h0;
      regVec_4010 <= 8'h0;
      regVec_4011 <= 8'h0;
      regVec_4012 <= 8'h0;
      regVec_4013 <= 8'h0;
      regVec_4014 <= 8'h0;
      regVec_4015 <= 8'h0;
      regVec_4016 <= 8'h0;
      regVec_4017 <= 8'h0;
      regVec_4018 <= 8'h0;
      regVec_4019 <= 8'h0;
      regVec_4020 <= 8'h0;
      regVec_4021 <= 8'h0;
      regVec_4022 <= 8'h0;
      regVec_4023 <= 8'h0;
      regVec_4024 <= 8'h0;
      regVec_4025 <= 8'h0;
      regVec_4026 <= 8'h0;
      regVec_4027 <= 8'h0;
      regVec_4028 <= 8'h0;
      regVec_4029 <= 8'h0;
      regVec_4030 <= 8'h0;
      regVec_4031 <= 8'h0;
      regVec_4032 <= 8'h0;
      regVec_4033 <= 8'h0;
      regVec_4034 <= 8'h0;
      regVec_4035 <= 8'h0;
      regVec_4036 <= 8'h0;
      regVec_4037 <= 8'h0;
      regVec_4038 <= 8'h0;
      regVec_4039 <= 8'h0;
      regVec_4040 <= 8'h0;
      regVec_4041 <= 8'h0;
      regVec_4042 <= 8'h0;
      regVec_4043 <= 8'h0;
      regVec_4044 <= 8'h0;
      regVec_4045 <= 8'h0;
      regVec_4046 <= 8'h0;
      regVec_4047 <= 8'h0;
      regVec_4048 <= 8'h0;
      regVec_4049 <= 8'h0;
      regVec_4050 <= 8'h0;
      regVec_4051 <= 8'h0;
      regVec_4052 <= 8'h0;
      regVec_4053 <= 8'h0;
      regVec_4054 <= 8'h0;
      regVec_4055 <= 8'h0;
      regVec_4056 <= 8'h0;
      regVec_4057 <= 8'h0;
      regVec_4058 <= 8'h0;
      regVec_4059 <= 8'h0;
      regVec_4060 <= 8'h0;
      regVec_4061 <= 8'h0;
      regVec_4062 <= 8'h0;
      regVec_4063 <= 8'h0;
      regVec_4064 <= 8'h0;
      regVec_4065 <= 8'h0;
      regVec_4066 <= 8'h0;
      regVec_4067 <= 8'h0;
      regVec_4068 <= 8'h0;
      regVec_4069 <= 8'h0;
      regVec_4070 <= 8'h0;
      regVec_4071 <= 8'h0;
      regVec_4072 <= 8'h0;
      regVec_4073 <= 8'h0;
      regVec_4074 <= 8'h0;
      regVec_4075 <= 8'h0;
      regVec_4076 <= 8'h0;
      regVec_4077 <= 8'h0;
      regVec_4078 <= 8'h0;
      regVec_4079 <= 8'h0;
      regVec_4080 <= 8'h0;
      regVec_4081 <= 8'h0;
      regVec_4082 <= 8'h0;
      regVec_4083 <= 8'h0;
      regVec_4084 <= 8'h0;
      regVec_4085 <= 8'h0;
      regVec_4086 <= 8'h0;
      regVec_4087 <= 8'h0;
      regVec_4088 <= 8'h0;
      regVec_4089 <= 8'h0;
      regVec_4090 <= 8'h0;
      regVec_4091 <= 8'h0;
      regVec_4092 <= 8'h0;
      regVec_4093 <= 8'h0;
      regVec_4094 <= 8'h0;
      regVec_4095 <= 8'h0;
      regAwAddr <= 12'h0;
      regAwId <= 4'b0000;
      regAwRegion <= 4'b0000;
      regAwLen <= 8'h0;
      regAwSize <= 3'b101;
      regAwBrust <= 2'b01;
      regAwLock <= 1'b0;
      regAwCache <= 4'b0000;
      regAwQos <= 4'b0000;
      regAwUser <= 1'b0;
      regAwProt <= 3'b000;
      regArAddr <= 12'h0;
      regArId <= 4'b0000;
      regArRegion <= 4'b0000;
      regArLen <= 8'h0;
      regArSize <= 3'b101;
      regArBrust <= 2'b01;
      regArLock <= 1'b0;
      regArCache <= 4'b0000;
      regArQos <= 4'b0000;
      regArUser <= 1'b0;
      regArProt <= 3'b000;
      updataAw <= 1'b1;
      writeSuccess <= 1'b0;
      updataAr <= 1'b1;
      rFireCounter_value <= 13'h0;
      AwArConflict <= 1'b0;
      regLast <= 1'b0;
    end else begin
      rFireCounter_value <= rFireCounter_valueNext;
      if(when_Axi4_transmission_l66) begin
        updataAw <= 1'b0;
      end else begin
        if(when_Axi4_transmission_l68) begin
          updataAw <= 1'b1;
        end
      end
      if(when_Axi4_transmission_l72) begin
        regAwAddr <= _zz_regAwAddr[11 : 0];
        regAwId <= axiSignal_aw_payload_id;
        regAwRegion <= axiSignal_aw_payload_region;
        regAwLen <= axiSignal_aw_payload_len;
        regAwSize <= axiSignal_aw_payload_size;
        regAwBrust <= axiSignal_aw_payload_burst;
        regAwLock <= axiSignal_aw_payload_lock;
        regAwCache <= axiSignal_aw_payload_cache;
        regAwQos <= axiSignal_aw_payload_qos;
        regAwUser <= axiSignal_aw_payload_user;
        regAwProt <= axiSignal_aw_payload_prot;
      end
      if(when_Axi4_transmission_l91) begin
        if(when_Axi4_transmission_l92) begin
          if(_zz_1[0]) begin
            regVec_0 <= _zz_regVec_0;
          end
          if(_zz_1[1]) begin
            regVec_1 <= _zz_regVec_0;
          end
          if(_zz_1[2]) begin
            regVec_2 <= _zz_regVec_0;
          end
          if(_zz_1[3]) begin
            regVec_3 <= _zz_regVec_0;
          end
          if(_zz_1[4]) begin
            regVec_4 <= _zz_regVec_0;
          end
          if(_zz_1[5]) begin
            regVec_5 <= _zz_regVec_0;
          end
          if(_zz_1[6]) begin
            regVec_6 <= _zz_regVec_0;
          end
          if(_zz_1[7]) begin
            regVec_7 <= _zz_regVec_0;
          end
          if(_zz_1[8]) begin
            regVec_8 <= _zz_regVec_0;
          end
          if(_zz_1[9]) begin
            regVec_9 <= _zz_regVec_0;
          end
          if(_zz_1[10]) begin
            regVec_10 <= _zz_regVec_0;
          end
          if(_zz_1[11]) begin
            regVec_11 <= _zz_regVec_0;
          end
          if(_zz_1[12]) begin
            regVec_12 <= _zz_regVec_0;
          end
          if(_zz_1[13]) begin
            regVec_13 <= _zz_regVec_0;
          end
          if(_zz_1[14]) begin
            regVec_14 <= _zz_regVec_0;
          end
          if(_zz_1[15]) begin
            regVec_15 <= _zz_regVec_0;
          end
          if(_zz_1[16]) begin
            regVec_16 <= _zz_regVec_0;
          end
          if(_zz_1[17]) begin
            regVec_17 <= _zz_regVec_0;
          end
          if(_zz_1[18]) begin
            regVec_18 <= _zz_regVec_0;
          end
          if(_zz_1[19]) begin
            regVec_19 <= _zz_regVec_0;
          end
          if(_zz_1[20]) begin
            regVec_20 <= _zz_regVec_0;
          end
          if(_zz_1[21]) begin
            regVec_21 <= _zz_regVec_0;
          end
          if(_zz_1[22]) begin
            regVec_22 <= _zz_regVec_0;
          end
          if(_zz_1[23]) begin
            regVec_23 <= _zz_regVec_0;
          end
          if(_zz_1[24]) begin
            regVec_24 <= _zz_regVec_0;
          end
          if(_zz_1[25]) begin
            regVec_25 <= _zz_regVec_0;
          end
          if(_zz_1[26]) begin
            regVec_26 <= _zz_regVec_0;
          end
          if(_zz_1[27]) begin
            regVec_27 <= _zz_regVec_0;
          end
          if(_zz_1[28]) begin
            regVec_28 <= _zz_regVec_0;
          end
          if(_zz_1[29]) begin
            regVec_29 <= _zz_regVec_0;
          end
          if(_zz_1[30]) begin
            regVec_30 <= _zz_regVec_0;
          end
          if(_zz_1[31]) begin
            regVec_31 <= _zz_regVec_0;
          end
          if(_zz_1[32]) begin
            regVec_32 <= _zz_regVec_0;
          end
          if(_zz_1[33]) begin
            regVec_33 <= _zz_regVec_0;
          end
          if(_zz_1[34]) begin
            regVec_34 <= _zz_regVec_0;
          end
          if(_zz_1[35]) begin
            regVec_35 <= _zz_regVec_0;
          end
          if(_zz_1[36]) begin
            regVec_36 <= _zz_regVec_0;
          end
          if(_zz_1[37]) begin
            regVec_37 <= _zz_regVec_0;
          end
          if(_zz_1[38]) begin
            regVec_38 <= _zz_regVec_0;
          end
          if(_zz_1[39]) begin
            regVec_39 <= _zz_regVec_0;
          end
          if(_zz_1[40]) begin
            regVec_40 <= _zz_regVec_0;
          end
          if(_zz_1[41]) begin
            regVec_41 <= _zz_regVec_0;
          end
          if(_zz_1[42]) begin
            regVec_42 <= _zz_regVec_0;
          end
          if(_zz_1[43]) begin
            regVec_43 <= _zz_regVec_0;
          end
          if(_zz_1[44]) begin
            regVec_44 <= _zz_regVec_0;
          end
          if(_zz_1[45]) begin
            regVec_45 <= _zz_regVec_0;
          end
          if(_zz_1[46]) begin
            regVec_46 <= _zz_regVec_0;
          end
          if(_zz_1[47]) begin
            regVec_47 <= _zz_regVec_0;
          end
          if(_zz_1[48]) begin
            regVec_48 <= _zz_regVec_0;
          end
          if(_zz_1[49]) begin
            regVec_49 <= _zz_regVec_0;
          end
          if(_zz_1[50]) begin
            regVec_50 <= _zz_regVec_0;
          end
          if(_zz_1[51]) begin
            regVec_51 <= _zz_regVec_0;
          end
          if(_zz_1[52]) begin
            regVec_52 <= _zz_regVec_0;
          end
          if(_zz_1[53]) begin
            regVec_53 <= _zz_regVec_0;
          end
          if(_zz_1[54]) begin
            regVec_54 <= _zz_regVec_0;
          end
          if(_zz_1[55]) begin
            regVec_55 <= _zz_regVec_0;
          end
          if(_zz_1[56]) begin
            regVec_56 <= _zz_regVec_0;
          end
          if(_zz_1[57]) begin
            regVec_57 <= _zz_regVec_0;
          end
          if(_zz_1[58]) begin
            regVec_58 <= _zz_regVec_0;
          end
          if(_zz_1[59]) begin
            regVec_59 <= _zz_regVec_0;
          end
          if(_zz_1[60]) begin
            regVec_60 <= _zz_regVec_0;
          end
          if(_zz_1[61]) begin
            regVec_61 <= _zz_regVec_0;
          end
          if(_zz_1[62]) begin
            regVec_62 <= _zz_regVec_0;
          end
          if(_zz_1[63]) begin
            regVec_63 <= _zz_regVec_0;
          end
          if(_zz_1[64]) begin
            regVec_64 <= _zz_regVec_0;
          end
          if(_zz_1[65]) begin
            regVec_65 <= _zz_regVec_0;
          end
          if(_zz_1[66]) begin
            regVec_66 <= _zz_regVec_0;
          end
          if(_zz_1[67]) begin
            regVec_67 <= _zz_regVec_0;
          end
          if(_zz_1[68]) begin
            regVec_68 <= _zz_regVec_0;
          end
          if(_zz_1[69]) begin
            regVec_69 <= _zz_regVec_0;
          end
          if(_zz_1[70]) begin
            regVec_70 <= _zz_regVec_0;
          end
          if(_zz_1[71]) begin
            regVec_71 <= _zz_regVec_0;
          end
          if(_zz_1[72]) begin
            regVec_72 <= _zz_regVec_0;
          end
          if(_zz_1[73]) begin
            regVec_73 <= _zz_regVec_0;
          end
          if(_zz_1[74]) begin
            regVec_74 <= _zz_regVec_0;
          end
          if(_zz_1[75]) begin
            regVec_75 <= _zz_regVec_0;
          end
          if(_zz_1[76]) begin
            regVec_76 <= _zz_regVec_0;
          end
          if(_zz_1[77]) begin
            regVec_77 <= _zz_regVec_0;
          end
          if(_zz_1[78]) begin
            regVec_78 <= _zz_regVec_0;
          end
          if(_zz_1[79]) begin
            regVec_79 <= _zz_regVec_0;
          end
          if(_zz_1[80]) begin
            regVec_80 <= _zz_regVec_0;
          end
          if(_zz_1[81]) begin
            regVec_81 <= _zz_regVec_0;
          end
          if(_zz_1[82]) begin
            regVec_82 <= _zz_regVec_0;
          end
          if(_zz_1[83]) begin
            regVec_83 <= _zz_regVec_0;
          end
          if(_zz_1[84]) begin
            regVec_84 <= _zz_regVec_0;
          end
          if(_zz_1[85]) begin
            regVec_85 <= _zz_regVec_0;
          end
          if(_zz_1[86]) begin
            regVec_86 <= _zz_regVec_0;
          end
          if(_zz_1[87]) begin
            regVec_87 <= _zz_regVec_0;
          end
          if(_zz_1[88]) begin
            regVec_88 <= _zz_regVec_0;
          end
          if(_zz_1[89]) begin
            regVec_89 <= _zz_regVec_0;
          end
          if(_zz_1[90]) begin
            regVec_90 <= _zz_regVec_0;
          end
          if(_zz_1[91]) begin
            regVec_91 <= _zz_regVec_0;
          end
          if(_zz_1[92]) begin
            regVec_92 <= _zz_regVec_0;
          end
          if(_zz_1[93]) begin
            regVec_93 <= _zz_regVec_0;
          end
          if(_zz_1[94]) begin
            regVec_94 <= _zz_regVec_0;
          end
          if(_zz_1[95]) begin
            regVec_95 <= _zz_regVec_0;
          end
          if(_zz_1[96]) begin
            regVec_96 <= _zz_regVec_0;
          end
          if(_zz_1[97]) begin
            regVec_97 <= _zz_regVec_0;
          end
          if(_zz_1[98]) begin
            regVec_98 <= _zz_regVec_0;
          end
          if(_zz_1[99]) begin
            regVec_99 <= _zz_regVec_0;
          end
          if(_zz_1[100]) begin
            regVec_100 <= _zz_regVec_0;
          end
          if(_zz_1[101]) begin
            regVec_101 <= _zz_regVec_0;
          end
          if(_zz_1[102]) begin
            regVec_102 <= _zz_regVec_0;
          end
          if(_zz_1[103]) begin
            regVec_103 <= _zz_regVec_0;
          end
          if(_zz_1[104]) begin
            regVec_104 <= _zz_regVec_0;
          end
          if(_zz_1[105]) begin
            regVec_105 <= _zz_regVec_0;
          end
          if(_zz_1[106]) begin
            regVec_106 <= _zz_regVec_0;
          end
          if(_zz_1[107]) begin
            regVec_107 <= _zz_regVec_0;
          end
          if(_zz_1[108]) begin
            regVec_108 <= _zz_regVec_0;
          end
          if(_zz_1[109]) begin
            regVec_109 <= _zz_regVec_0;
          end
          if(_zz_1[110]) begin
            regVec_110 <= _zz_regVec_0;
          end
          if(_zz_1[111]) begin
            regVec_111 <= _zz_regVec_0;
          end
          if(_zz_1[112]) begin
            regVec_112 <= _zz_regVec_0;
          end
          if(_zz_1[113]) begin
            regVec_113 <= _zz_regVec_0;
          end
          if(_zz_1[114]) begin
            regVec_114 <= _zz_regVec_0;
          end
          if(_zz_1[115]) begin
            regVec_115 <= _zz_regVec_0;
          end
          if(_zz_1[116]) begin
            regVec_116 <= _zz_regVec_0;
          end
          if(_zz_1[117]) begin
            regVec_117 <= _zz_regVec_0;
          end
          if(_zz_1[118]) begin
            regVec_118 <= _zz_regVec_0;
          end
          if(_zz_1[119]) begin
            regVec_119 <= _zz_regVec_0;
          end
          if(_zz_1[120]) begin
            regVec_120 <= _zz_regVec_0;
          end
          if(_zz_1[121]) begin
            regVec_121 <= _zz_regVec_0;
          end
          if(_zz_1[122]) begin
            regVec_122 <= _zz_regVec_0;
          end
          if(_zz_1[123]) begin
            regVec_123 <= _zz_regVec_0;
          end
          if(_zz_1[124]) begin
            regVec_124 <= _zz_regVec_0;
          end
          if(_zz_1[125]) begin
            regVec_125 <= _zz_regVec_0;
          end
          if(_zz_1[126]) begin
            regVec_126 <= _zz_regVec_0;
          end
          if(_zz_1[127]) begin
            regVec_127 <= _zz_regVec_0;
          end
          if(_zz_1[128]) begin
            regVec_128 <= _zz_regVec_0;
          end
          if(_zz_1[129]) begin
            regVec_129 <= _zz_regVec_0;
          end
          if(_zz_1[130]) begin
            regVec_130 <= _zz_regVec_0;
          end
          if(_zz_1[131]) begin
            regVec_131 <= _zz_regVec_0;
          end
          if(_zz_1[132]) begin
            regVec_132 <= _zz_regVec_0;
          end
          if(_zz_1[133]) begin
            regVec_133 <= _zz_regVec_0;
          end
          if(_zz_1[134]) begin
            regVec_134 <= _zz_regVec_0;
          end
          if(_zz_1[135]) begin
            regVec_135 <= _zz_regVec_0;
          end
          if(_zz_1[136]) begin
            regVec_136 <= _zz_regVec_0;
          end
          if(_zz_1[137]) begin
            regVec_137 <= _zz_regVec_0;
          end
          if(_zz_1[138]) begin
            regVec_138 <= _zz_regVec_0;
          end
          if(_zz_1[139]) begin
            regVec_139 <= _zz_regVec_0;
          end
          if(_zz_1[140]) begin
            regVec_140 <= _zz_regVec_0;
          end
          if(_zz_1[141]) begin
            regVec_141 <= _zz_regVec_0;
          end
          if(_zz_1[142]) begin
            regVec_142 <= _zz_regVec_0;
          end
          if(_zz_1[143]) begin
            regVec_143 <= _zz_regVec_0;
          end
          if(_zz_1[144]) begin
            regVec_144 <= _zz_regVec_0;
          end
          if(_zz_1[145]) begin
            regVec_145 <= _zz_regVec_0;
          end
          if(_zz_1[146]) begin
            regVec_146 <= _zz_regVec_0;
          end
          if(_zz_1[147]) begin
            regVec_147 <= _zz_regVec_0;
          end
          if(_zz_1[148]) begin
            regVec_148 <= _zz_regVec_0;
          end
          if(_zz_1[149]) begin
            regVec_149 <= _zz_regVec_0;
          end
          if(_zz_1[150]) begin
            regVec_150 <= _zz_regVec_0;
          end
          if(_zz_1[151]) begin
            regVec_151 <= _zz_regVec_0;
          end
          if(_zz_1[152]) begin
            regVec_152 <= _zz_regVec_0;
          end
          if(_zz_1[153]) begin
            regVec_153 <= _zz_regVec_0;
          end
          if(_zz_1[154]) begin
            regVec_154 <= _zz_regVec_0;
          end
          if(_zz_1[155]) begin
            regVec_155 <= _zz_regVec_0;
          end
          if(_zz_1[156]) begin
            regVec_156 <= _zz_regVec_0;
          end
          if(_zz_1[157]) begin
            regVec_157 <= _zz_regVec_0;
          end
          if(_zz_1[158]) begin
            regVec_158 <= _zz_regVec_0;
          end
          if(_zz_1[159]) begin
            regVec_159 <= _zz_regVec_0;
          end
          if(_zz_1[160]) begin
            regVec_160 <= _zz_regVec_0;
          end
          if(_zz_1[161]) begin
            regVec_161 <= _zz_regVec_0;
          end
          if(_zz_1[162]) begin
            regVec_162 <= _zz_regVec_0;
          end
          if(_zz_1[163]) begin
            regVec_163 <= _zz_regVec_0;
          end
          if(_zz_1[164]) begin
            regVec_164 <= _zz_regVec_0;
          end
          if(_zz_1[165]) begin
            regVec_165 <= _zz_regVec_0;
          end
          if(_zz_1[166]) begin
            regVec_166 <= _zz_regVec_0;
          end
          if(_zz_1[167]) begin
            regVec_167 <= _zz_regVec_0;
          end
          if(_zz_1[168]) begin
            regVec_168 <= _zz_regVec_0;
          end
          if(_zz_1[169]) begin
            regVec_169 <= _zz_regVec_0;
          end
          if(_zz_1[170]) begin
            regVec_170 <= _zz_regVec_0;
          end
          if(_zz_1[171]) begin
            regVec_171 <= _zz_regVec_0;
          end
          if(_zz_1[172]) begin
            regVec_172 <= _zz_regVec_0;
          end
          if(_zz_1[173]) begin
            regVec_173 <= _zz_regVec_0;
          end
          if(_zz_1[174]) begin
            regVec_174 <= _zz_regVec_0;
          end
          if(_zz_1[175]) begin
            regVec_175 <= _zz_regVec_0;
          end
          if(_zz_1[176]) begin
            regVec_176 <= _zz_regVec_0;
          end
          if(_zz_1[177]) begin
            regVec_177 <= _zz_regVec_0;
          end
          if(_zz_1[178]) begin
            regVec_178 <= _zz_regVec_0;
          end
          if(_zz_1[179]) begin
            regVec_179 <= _zz_regVec_0;
          end
          if(_zz_1[180]) begin
            regVec_180 <= _zz_regVec_0;
          end
          if(_zz_1[181]) begin
            regVec_181 <= _zz_regVec_0;
          end
          if(_zz_1[182]) begin
            regVec_182 <= _zz_regVec_0;
          end
          if(_zz_1[183]) begin
            regVec_183 <= _zz_regVec_0;
          end
          if(_zz_1[184]) begin
            regVec_184 <= _zz_regVec_0;
          end
          if(_zz_1[185]) begin
            regVec_185 <= _zz_regVec_0;
          end
          if(_zz_1[186]) begin
            regVec_186 <= _zz_regVec_0;
          end
          if(_zz_1[187]) begin
            regVec_187 <= _zz_regVec_0;
          end
          if(_zz_1[188]) begin
            regVec_188 <= _zz_regVec_0;
          end
          if(_zz_1[189]) begin
            regVec_189 <= _zz_regVec_0;
          end
          if(_zz_1[190]) begin
            regVec_190 <= _zz_regVec_0;
          end
          if(_zz_1[191]) begin
            regVec_191 <= _zz_regVec_0;
          end
          if(_zz_1[192]) begin
            regVec_192 <= _zz_regVec_0;
          end
          if(_zz_1[193]) begin
            regVec_193 <= _zz_regVec_0;
          end
          if(_zz_1[194]) begin
            regVec_194 <= _zz_regVec_0;
          end
          if(_zz_1[195]) begin
            regVec_195 <= _zz_regVec_0;
          end
          if(_zz_1[196]) begin
            regVec_196 <= _zz_regVec_0;
          end
          if(_zz_1[197]) begin
            regVec_197 <= _zz_regVec_0;
          end
          if(_zz_1[198]) begin
            regVec_198 <= _zz_regVec_0;
          end
          if(_zz_1[199]) begin
            regVec_199 <= _zz_regVec_0;
          end
          if(_zz_1[200]) begin
            regVec_200 <= _zz_regVec_0;
          end
          if(_zz_1[201]) begin
            regVec_201 <= _zz_regVec_0;
          end
          if(_zz_1[202]) begin
            regVec_202 <= _zz_regVec_0;
          end
          if(_zz_1[203]) begin
            regVec_203 <= _zz_regVec_0;
          end
          if(_zz_1[204]) begin
            regVec_204 <= _zz_regVec_0;
          end
          if(_zz_1[205]) begin
            regVec_205 <= _zz_regVec_0;
          end
          if(_zz_1[206]) begin
            regVec_206 <= _zz_regVec_0;
          end
          if(_zz_1[207]) begin
            regVec_207 <= _zz_regVec_0;
          end
          if(_zz_1[208]) begin
            regVec_208 <= _zz_regVec_0;
          end
          if(_zz_1[209]) begin
            regVec_209 <= _zz_regVec_0;
          end
          if(_zz_1[210]) begin
            regVec_210 <= _zz_regVec_0;
          end
          if(_zz_1[211]) begin
            regVec_211 <= _zz_regVec_0;
          end
          if(_zz_1[212]) begin
            regVec_212 <= _zz_regVec_0;
          end
          if(_zz_1[213]) begin
            regVec_213 <= _zz_regVec_0;
          end
          if(_zz_1[214]) begin
            regVec_214 <= _zz_regVec_0;
          end
          if(_zz_1[215]) begin
            regVec_215 <= _zz_regVec_0;
          end
          if(_zz_1[216]) begin
            regVec_216 <= _zz_regVec_0;
          end
          if(_zz_1[217]) begin
            regVec_217 <= _zz_regVec_0;
          end
          if(_zz_1[218]) begin
            regVec_218 <= _zz_regVec_0;
          end
          if(_zz_1[219]) begin
            regVec_219 <= _zz_regVec_0;
          end
          if(_zz_1[220]) begin
            regVec_220 <= _zz_regVec_0;
          end
          if(_zz_1[221]) begin
            regVec_221 <= _zz_regVec_0;
          end
          if(_zz_1[222]) begin
            regVec_222 <= _zz_regVec_0;
          end
          if(_zz_1[223]) begin
            regVec_223 <= _zz_regVec_0;
          end
          if(_zz_1[224]) begin
            regVec_224 <= _zz_regVec_0;
          end
          if(_zz_1[225]) begin
            regVec_225 <= _zz_regVec_0;
          end
          if(_zz_1[226]) begin
            regVec_226 <= _zz_regVec_0;
          end
          if(_zz_1[227]) begin
            regVec_227 <= _zz_regVec_0;
          end
          if(_zz_1[228]) begin
            regVec_228 <= _zz_regVec_0;
          end
          if(_zz_1[229]) begin
            regVec_229 <= _zz_regVec_0;
          end
          if(_zz_1[230]) begin
            regVec_230 <= _zz_regVec_0;
          end
          if(_zz_1[231]) begin
            regVec_231 <= _zz_regVec_0;
          end
          if(_zz_1[232]) begin
            regVec_232 <= _zz_regVec_0;
          end
          if(_zz_1[233]) begin
            regVec_233 <= _zz_regVec_0;
          end
          if(_zz_1[234]) begin
            regVec_234 <= _zz_regVec_0;
          end
          if(_zz_1[235]) begin
            regVec_235 <= _zz_regVec_0;
          end
          if(_zz_1[236]) begin
            regVec_236 <= _zz_regVec_0;
          end
          if(_zz_1[237]) begin
            regVec_237 <= _zz_regVec_0;
          end
          if(_zz_1[238]) begin
            regVec_238 <= _zz_regVec_0;
          end
          if(_zz_1[239]) begin
            regVec_239 <= _zz_regVec_0;
          end
          if(_zz_1[240]) begin
            regVec_240 <= _zz_regVec_0;
          end
          if(_zz_1[241]) begin
            regVec_241 <= _zz_regVec_0;
          end
          if(_zz_1[242]) begin
            regVec_242 <= _zz_regVec_0;
          end
          if(_zz_1[243]) begin
            regVec_243 <= _zz_regVec_0;
          end
          if(_zz_1[244]) begin
            regVec_244 <= _zz_regVec_0;
          end
          if(_zz_1[245]) begin
            regVec_245 <= _zz_regVec_0;
          end
          if(_zz_1[246]) begin
            regVec_246 <= _zz_regVec_0;
          end
          if(_zz_1[247]) begin
            regVec_247 <= _zz_regVec_0;
          end
          if(_zz_1[248]) begin
            regVec_248 <= _zz_regVec_0;
          end
          if(_zz_1[249]) begin
            regVec_249 <= _zz_regVec_0;
          end
          if(_zz_1[250]) begin
            regVec_250 <= _zz_regVec_0;
          end
          if(_zz_1[251]) begin
            regVec_251 <= _zz_regVec_0;
          end
          if(_zz_1[252]) begin
            regVec_252 <= _zz_regVec_0;
          end
          if(_zz_1[253]) begin
            regVec_253 <= _zz_regVec_0;
          end
          if(_zz_1[254]) begin
            regVec_254 <= _zz_regVec_0;
          end
          if(_zz_1[255]) begin
            regVec_255 <= _zz_regVec_0;
          end
          if(_zz_1[256]) begin
            regVec_256 <= _zz_regVec_0;
          end
          if(_zz_1[257]) begin
            regVec_257 <= _zz_regVec_0;
          end
          if(_zz_1[258]) begin
            regVec_258 <= _zz_regVec_0;
          end
          if(_zz_1[259]) begin
            regVec_259 <= _zz_regVec_0;
          end
          if(_zz_1[260]) begin
            regVec_260 <= _zz_regVec_0;
          end
          if(_zz_1[261]) begin
            regVec_261 <= _zz_regVec_0;
          end
          if(_zz_1[262]) begin
            regVec_262 <= _zz_regVec_0;
          end
          if(_zz_1[263]) begin
            regVec_263 <= _zz_regVec_0;
          end
          if(_zz_1[264]) begin
            regVec_264 <= _zz_regVec_0;
          end
          if(_zz_1[265]) begin
            regVec_265 <= _zz_regVec_0;
          end
          if(_zz_1[266]) begin
            regVec_266 <= _zz_regVec_0;
          end
          if(_zz_1[267]) begin
            regVec_267 <= _zz_regVec_0;
          end
          if(_zz_1[268]) begin
            regVec_268 <= _zz_regVec_0;
          end
          if(_zz_1[269]) begin
            regVec_269 <= _zz_regVec_0;
          end
          if(_zz_1[270]) begin
            regVec_270 <= _zz_regVec_0;
          end
          if(_zz_1[271]) begin
            regVec_271 <= _zz_regVec_0;
          end
          if(_zz_1[272]) begin
            regVec_272 <= _zz_regVec_0;
          end
          if(_zz_1[273]) begin
            regVec_273 <= _zz_regVec_0;
          end
          if(_zz_1[274]) begin
            regVec_274 <= _zz_regVec_0;
          end
          if(_zz_1[275]) begin
            regVec_275 <= _zz_regVec_0;
          end
          if(_zz_1[276]) begin
            regVec_276 <= _zz_regVec_0;
          end
          if(_zz_1[277]) begin
            regVec_277 <= _zz_regVec_0;
          end
          if(_zz_1[278]) begin
            regVec_278 <= _zz_regVec_0;
          end
          if(_zz_1[279]) begin
            regVec_279 <= _zz_regVec_0;
          end
          if(_zz_1[280]) begin
            regVec_280 <= _zz_regVec_0;
          end
          if(_zz_1[281]) begin
            regVec_281 <= _zz_regVec_0;
          end
          if(_zz_1[282]) begin
            regVec_282 <= _zz_regVec_0;
          end
          if(_zz_1[283]) begin
            regVec_283 <= _zz_regVec_0;
          end
          if(_zz_1[284]) begin
            regVec_284 <= _zz_regVec_0;
          end
          if(_zz_1[285]) begin
            regVec_285 <= _zz_regVec_0;
          end
          if(_zz_1[286]) begin
            regVec_286 <= _zz_regVec_0;
          end
          if(_zz_1[287]) begin
            regVec_287 <= _zz_regVec_0;
          end
          if(_zz_1[288]) begin
            regVec_288 <= _zz_regVec_0;
          end
          if(_zz_1[289]) begin
            regVec_289 <= _zz_regVec_0;
          end
          if(_zz_1[290]) begin
            regVec_290 <= _zz_regVec_0;
          end
          if(_zz_1[291]) begin
            regVec_291 <= _zz_regVec_0;
          end
          if(_zz_1[292]) begin
            regVec_292 <= _zz_regVec_0;
          end
          if(_zz_1[293]) begin
            regVec_293 <= _zz_regVec_0;
          end
          if(_zz_1[294]) begin
            regVec_294 <= _zz_regVec_0;
          end
          if(_zz_1[295]) begin
            regVec_295 <= _zz_regVec_0;
          end
          if(_zz_1[296]) begin
            regVec_296 <= _zz_regVec_0;
          end
          if(_zz_1[297]) begin
            regVec_297 <= _zz_regVec_0;
          end
          if(_zz_1[298]) begin
            regVec_298 <= _zz_regVec_0;
          end
          if(_zz_1[299]) begin
            regVec_299 <= _zz_regVec_0;
          end
          if(_zz_1[300]) begin
            regVec_300 <= _zz_regVec_0;
          end
          if(_zz_1[301]) begin
            regVec_301 <= _zz_regVec_0;
          end
          if(_zz_1[302]) begin
            regVec_302 <= _zz_regVec_0;
          end
          if(_zz_1[303]) begin
            regVec_303 <= _zz_regVec_0;
          end
          if(_zz_1[304]) begin
            regVec_304 <= _zz_regVec_0;
          end
          if(_zz_1[305]) begin
            regVec_305 <= _zz_regVec_0;
          end
          if(_zz_1[306]) begin
            regVec_306 <= _zz_regVec_0;
          end
          if(_zz_1[307]) begin
            regVec_307 <= _zz_regVec_0;
          end
          if(_zz_1[308]) begin
            regVec_308 <= _zz_regVec_0;
          end
          if(_zz_1[309]) begin
            regVec_309 <= _zz_regVec_0;
          end
          if(_zz_1[310]) begin
            regVec_310 <= _zz_regVec_0;
          end
          if(_zz_1[311]) begin
            regVec_311 <= _zz_regVec_0;
          end
          if(_zz_1[312]) begin
            regVec_312 <= _zz_regVec_0;
          end
          if(_zz_1[313]) begin
            regVec_313 <= _zz_regVec_0;
          end
          if(_zz_1[314]) begin
            regVec_314 <= _zz_regVec_0;
          end
          if(_zz_1[315]) begin
            regVec_315 <= _zz_regVec_0;
          end
          if(_zz_1[316]) begin
            regVec_316 <= _zz_regVec_0;
          end
          if(_zz_1[317]) begin
            regVec_317 <= _zz_regVec_0;
          end
          if(_zz_1[318]) begin
            regVec_318 <= _zz_regVec_0;
          end
          if(_zz_1[319]) begin
            regVec_319 <= _zz_regVec_0;
          end
          if(_zz_1[320]) begin
            regVec_320 <= _zz_regVec_0;
          end
          if(_zz_1[321]) begin
            regVec_321 <= _zz_regVec_0;
          end
          if(_zz_1[322]) begin
            regVec_322 <= _zz_regVec_0;
          end
          if(_zz_1[323]) begin
            regVec_323 <= _zz_regVec_0;
          end
          if(_zz_1[324]) begin
            regVec_324 <= _zz_regVec_0;
          end
          if(_zz_1[325]) begin
            regVec_325 <= _zz_regVec_0;
          end
          if(_zz_1[326]) begin
            regVec_326 <= _zz_regVec_0;
          end
          if(_zz_1[327]) begin
            regVec_327 <= _zz_regVec_0;
          end
          if(_zz_1[328]) begin
            regVec_328 <= _zz_regVec_0;
          end
          if(_zz_1[329]) begin
            regVec_329 <= _zz_regVec_0;
          end
          if(_zz_1[330]) begin
            regVec_330 <= _zz_regVec_0;
          end
          if(_zz_1[331]) begin
            regVec_331 <= _zz_regVec_0;
          end
          if(_zz_1[332]) begin
            regVec_332 <= _zz_regVec_0;
          end
          if(_zz_1[333]) begin
            regVec_333 <= _zz_regVec_0;
          end
          if(_zz_1[334]) begin
            regVec_334 <= _zz_regVec_0;
          end
          if(_zz_1[335]) begin
            regVec_335 <= _zz_regVec_0;
          end
          if(_zz_1[336]) begin
            regVec_336 <= _zz_regVec_0;
          end
          if(_zz_1[337]) begin
            regVec_337 <= _zz_regVec_0;
          end
          if(_zz_1[338]) begin
            regVec_338 <= _zz_regVec_0;
          end
          if(_zz_1[339]) begin
            regVec_339 <= _zz_regVec_0;
          end
          if(_zz_1[340]) begin
            regVec_340 <= _zz_regVec_0;
          end
          if(_zz_1[341]) begin
            regVec_341 <= _zz_regVec_0;
          end
          if(_zz_1[342]) begin
            regVec_342 <= _zz_regVec_0;
          end
          if(_zz_1[343]) begin
            regVec_343 <= _zz_regVec_0;
          end
          if(_zz_1[344]) begin
            regVec_344 <= _zz_regVec_0;
          end
          if(_zz_1[345]) begin
            regVec_345 <= _zz_regVec_0;
          end
          if(_zz_1[346]) begin
            regVec_346 <= _zz_regVec_0;
          end
          if(_zz_1[347]) begin
            regVec_347 <= _zz_regVec_0;
          end
          if(_zz_1[348]) begin
            regVec_348 <= _zz_regVec_0;
          end
          if(_zz_1[349]) begin
            regVec_349 <= _zz_regVec_0;
          end
          if(_zz_1[350]) begin
            regVec_350 <= _zz_regVec_0;
          end
          if(_zz_1[351]) begin
            regVec_351 <= _zz_regVec_0;
          end
          if(_zz_1[352]) begin
            regVec_352 <= _zz_regVec_0;
          end
          if(_zz_1[353]) begin
            regVec_353 <= _zz_regVec_0;
          end
          if(_zz_1[354]) begin
            regVec_354 <= _zz_regVec_0;
          end
          if(_zz_1[355]) begin
            regVec_355 <= _zz_regVec_0;
          end
          if(_zz_1[356]) begin
            regVec_356 <= _zz_regVec_0;
          end
          if(_zz_1[357]) begin
            regVec_357 <= _zz_regVec_0;
          end
          if(_zz_1[358]) begin
            regVec_358 <= _zz_regVec_0;
          end
          if(_zz_1[359]) begin
            regVec_359 <= _zz_regVec_0;
          end
          if(_zz_1[360]) begin
            regVec_360 <= _zz_regVec_0;
          end
          if(_zz_1[361]) begin
            regVec_361 <= _zz_regVec_0;
          end
          if(_zz_1[362]) begin
            regVec_362 <= _zz_regVec_0;
          end
          if(_zz_1[363]) begin
            regVec_363 <= _zz_regVec_0;
          end
          if(_zz_1[364]) begin
            regVec_364 <= _zz_regVec_0;
          end
          if(_zz_1[365]) begin
            regVec_365 <= _zz_regVec_0;
          end
          if(_zz_1[366]) begin
            regVec_366 <= _zz_regVec_0;
          end
          if(_zz_1[367]) begin
            regVec_367 <= _zz_regVec_0;
          end
          if(_zz_1[368]) begin
            regVec_368 <= _zz_regVec_0;
          end
          if(_zz_1[369]) begin
            regVec_369 <= _zz_regVec_0;
          end
          if(_zz_1[370]) begin
            regVec_370 <= _zz_regVec_0;
          end
          if(_zz_1[371]) begin
            regVec_371 <= _zz_regVec_0;
          end
          if(_zz_1[372]) begin
            regVec_372 <= _zz_regVec_0;
          end
          if(_zz_1[373]) begin
            regVec_373 <= _zz_regVec_0;
          end
          if(_zz_1[374]) begin
            regVec_374 <= _zz_regVec_0;
          end
          if(_zz_1[375]) begin
            regVec_375 <= _zz_regVec_0;
          end
          if(_zz_1[376]) begin
            regVec_376 <= _zz_regVec_0;
          end
          if(_zz_1[377]) begin
            regVec_377 <= _zz_regVec_0;
          end
          if(_zz_1[378]) begin
            regVec_378 <= _zz_regVec_0;
          end
          if(_zz_1[379]) begin
            regVec_379 <= _zz_regVec_0;
          end
          if(_zz_1[380]) begin
            regVec_380 <= _zz_regVec_0;
          end
          if(_zz_1[381]) begin
            regVec_381 <= _zz_regVec_0;
          end
          if(_zz_1[382]) begin
            regVec_382 <= _zz_regVec_0;
          end
          if(_zz_1[383]) begin
            regVec_383 <= _zz_regVec_0;
          end
          if(_zz_1[384]) begin
            regVec_384 <= _zz_regVec_0;
          end
          if(_zz_1[385]) begin
            regVec_385 <= _zz_regVec_0;
          end
          if(_zz_1[386]) begin
            regVec_386 <= _zz_regVec_0;
          end
          if(_zz_1[387]) begin
            regVec_387 <= _zz_regVec_0;
          end
          if(_zz_1[388]) begin
            regVec_388 <= _zz_regVec_0;
          end
          if(_zz_1[389]) begin
            regVec_389 <= _zz_regVec_0;
          end
          if(_zz_1[390]) begin
            regVec_390 <= _zz_regVec_0;
          end
          if(_zz_1[391]) begin
            regVec_391 <= _zz_regVec_0;
          end
          if(_zz_1[392]) begin
            regVec_392 <= _zz_regVec_0;
          end
          if(_zz_1[393]) begin
            regVec_393 <= _zz_regVec_0;
          end
          if(_zz_1[394]) begin
            regVec_394 <= _zz_regVec_0;
          end
          if(_zz_1[395]) begin
            regVec_395 <= _zz_regVec_0;
          end
          if(_zz_1[396]) begin
            regVec_396 <= _zz_regVec_0;
          end
          if(_zz_1[397]) begin
            regVec_397 <= _zz_regVec_0;
          end
          if(_zz_1[398]) begin
            regVec_398 <= _zz_regVec_0;
          end
          if(_zz_1[399]) begin
            regVec_399 <= _zz_regVec_0;
          end
          if(_zz_1[400]) begin
            regVec_400 <= _zz_regVec_0;
          end
          if(_zz_1[401]) begin
            regVec_401 <= _zz_regVec_0;
          end
          if(_zz_1[402]) begin
            regVec_402 <= _zz_regVec_0;
          end
          if(_zz_1[403]) begin
            regVec_403 <= _zz_regVec_0;
          end
          if(_zz_1[404]) begin
            regVec_404 <= _zz_regVec_0;
          end
          if(_zz_1[405]) begin
            regVec_405 <= _zz_regVec_0;
          end
          if(_zz_1[406]) begin
            regVec_406 <= _zz_regVec_0;
          end
          if(_zz_1[407]) begin
            regVec_407 <= _zz_regVec_0;
          end
          if(_zz_1[408]) begin
            regVec_408 <= _zz_regVec_0;
          end
          if(_zz_1[409]) begin
            regVec_409 <= _zz_regVec_0;
          end
          if(_zz_1[410]) begin
            regVec_410 <= _zz_regVec_0;
          end
          if(_zz_1[411]) begin
            regVec_411 <= _zz_regVec_0;
          end
          if(_zz_1[412]) begin
            regVec_412 <= _zz_regVec_0;
          end
          if(_zz_1[413]) begin
            regVec_413 <= _zz_regVec_0;
          end
          if(_zz_1[414]) begin
            regVec_414 <= _zz_regVec_0;
          end
          if(_zz_1[415]) begin
            regVec_415 <= _zz_regVec_0;
          end
          if(_zz_1[416]) begin
            regVec_416 <= _zz_regVec_0;
          end
          if(_zz_1[417]) begin
            regVec_417 <= _zz_regVec_0;
          end
          if(_zz_1[418]) begin
            regVec_418 <= _zz_regVec_0;
          end
          if(_zz_1[419]) begin
            regVec_419 <= _zz_regVec_0;
          end
          if(_zz_1[420]) begin
            regVec_420 <= _zz_regVec_0;
          end
          if(_zz_1[421]) begin
            regVec_421 <= _zz_regVec_0;
          end
          if(_zz_1[422]) begin
            regVec_422 <= _zz_regVec_0;
          end
          if(_zz_1[423]) begin
            regVec_423 <= _zz_regVec_0;
          end
          if(_zz_1[424]) begin
            regVec_424 <= _zz_regVec_0;
          end
          if(_zz_1[425]) begin
            regVec_425 <= _zz_regVec_0;
          end
          if(_zz_1[426]) begin
            regVec_426 <= _zz_regVec_0;
          end
          if(_zz_1[427]) begin
            regVec_427 <= _zz_regVec_0;
          end
          if(_zz_1[428]) begin
            regVec_428 <= _zz_regVec_0;
          end
          if(_zz_1[429]) begin
            regVec_429 <= _zz_regVec_0;
          end
          if(_zz_1[430]) begin
            regVec_430 <= _zz_regVec_0;
          end
          if(_zz_1[431]) begin
            regVec_431 <= _zz_regVec_0;
          end
          if(_zz_1[432]) begin
            regVec_432 <= _zz_regVec_0;
          end
          if(_zz_1[433]) begin
            regVec_433 <= _zz_regVec_0;
          end
          if(_zz_1[434]) begin
            regVec_434 <= _zz_regVec_0;
          end
          if(_zz_1[435]) begin
            regVec_435 <= _zz_regVec_0;
          end
          if(_zz_1[436]) begin
            regVec_436 <= _zz_regVec_0;
          end
          if(_zz_1[437]) begin
            regVec_437 <= _zz_regVec_0;
          end
          if(_zz_1[438]) begin
            regVec_438 <= _zz_regVec_0;
          end
          if(_zz_1[439]) begin
            regVec_439 <= _zz_regVec_0;
          end
          if(_zz_1[440]) begin
            regVec_440 <= _zz_regVec_0;
          end
          if(_zz_1[441]) begin
            regVec_441 <= _zz_regVec_0;
          end
          if(_zz_1[442]) begin
            regVec_442 <= _zz_regVec_0;
          end
          if(_zz_1[443]) begin
            regVec_443 <= _zz_regVec_0;
          end
          if(_zz_1[444]) begin
            regVec_444 <= _zz_regVec_0;
          end
          if(_zz_1[445]) begin
            regVec_445 <= _zz_regVec_0;
          end
          if(_zz_1[446]) begin
            regVec_446 <= _zz_regVec_0;
          end
          if(_zz_1[447]) begin
            regVec_447 <= _zz_regVec_0;
          end
          if(_zz_1[448]) begin
            regVec_448 <= _zz_regVec_0;
          end
          if(_zz_1[449]) begin
            regVec_449 <= _zz_regVec_0;
          end
          if(_zz_1[450]) begin
            regVec_450 <= _zz_regVec_0;
          end
          if(_zz_1[451]) begin
            regVec_451 <= _zz_regVec_0;
          end
          if(_zz_1[452]) begin
            regVec_452 <= _zz_regVec_0;
          end
          if(_zz_1[453]) begin
            regVec_453 <= _zz_regVec_0;
          end
          if(_zz_1[454]) begin
            regVec_454 <= _zz_regVec_0;
          end
          if(_zz_1[455]) begin
            regVec_455 <= _zz_regVec_0;
          end
          if(_zz_1[456]) begin
            regVec_456 <= _zz_regVec_0;
          end
          if(_zz_1[457]) begin
            regVec_457 <= _zz_regVec_0;
          end
          if(_zz_1[458]) begin
            regVec_458 <= _zz_regVec_0;
          end
          if(_zz_1[459]) begin
            regVec_459 <= _zz_regVec_0;
          end
          if(_zz_1[460]) begin
            regVec_460 <= _zz_regVec_0;
          end
          if(_zz_1[461]) begin
            regVec_461 <= _zz_regVec_0;
          end
          if(_zz_1[462]) begin
            regVec_462 <= _zz_regVec_0;
          end
          if(_zz_1[463]) begin
            regVec_463 <= _zz_regVec_0;
          end
          if(_zz_1[464]) begin
            regVec_464 <= _zz_regVec_0;
          end
          if(_zz_1[465]) begin
            regVec_465 <= _zz_regVec_0;
          end
          if(_zz_1[466]) begin
            regVec_466 <= _zz_regVec_0;
          end
          if(_zz_1[467]) begin
            regVec_467 <= _zz_regVec_0;
          end
          if(_zz_1[468]) begin
            regVec_468 <= _zz_regVec_0;
          end
          if(_zz_1[469]) begin
            regVec_469 <= _zz_regVec_0;
          end
          if(_zz_1[470]) begin
            regVec_470 <= _zz_regVec_0;
          end
          if(_zz_1[471]) begin
            regVec_471 <= _zz_regVec_0;
          end
          if(_zz_1[472]) begin
            regVec_472 <= _zz_regVec_0;
          end
          if(_zz_1[473]) begin
            regVec_473 <= _zz_regVec_0;
          end
          if(_zz_1[474]) begin
            regVec_474 <= _zz_regVec_0;
          end
          if(_zz_1[475]) begin
            regVec_475 <= _zz_regVec_0;
          end
          if(_zz_1[476]) begin
            regVec_476 <= _zz_regVec_0;
          end
          if(_zz_1[477]) begin
            regVec_477 <= _zz_regVec_0;
          end
          if(_zz_1[478]) begin
            regVec_478 <= _zz_regVec_0;
          end
          if(_zz_1[479]) begin
            regVec_479 <= _zz_regVec_0;
          end
          if(_zz_1[480]) begin
            regVec_480 <= _zz_regVec_0;
          end
          if(_zz_1[481]) begin
            regVec_481 <= _zz_regVec_0;
          end
          if(_zz_1[482]) begin
            regVec_482 <= _zz_regVec_0;
          end
          if(_zz_1[483]) begin
            regVec_483 <= _zz_regVec_0;
          end
          if(_zz_1[484]) begin
            regVec_484 <= _zz_regVec_0;
          end
          if(_zz_1[485]) begin
            regVec_485 <= _zz_regVec_0;
          end
          if(_zz_1[486]) begin
            regVec_486 <= _zz_regVec_0;
          end
          if(_zz_1[487]) begin
            regVec_487 <= _zz_regVec_0;
          end
          if(_zz_1[488]) begin
            regVec_488 <= _zz_regVec_0;
          end
          if(_zz_1[489]) begin
            regVec_489 <= _zz_regVec_0;
          end
          if(_zz_1[490]) begin
            regVec_490 <= _zz_regVec_0;
          end
          if(_zz_1[491]) begin
            regVec_491 <= _zz_regVec_0;
          end
          if(_zz_1[492]) begin
            regVec_492 <= _zz_regVec_0;
          end
          if(_zz_1[493]) begin
            regVec_493 <= _zz_regVec_0;
          end
          if(_zz_1[494]) begin
            regVec_494 <= _zz_regVec_0;
          end
          if(_zz_1[495]) begin
            regVec_495 <= _zz_regVec_0;
          end
          if(_zz_1[496]) begin
            regVec_496 <= _zz_regVec_0;
          end
          if(_zz_1[497]) begin
            regVec_497 <= _zz_regVec_0;
          end
          if(_zz_1[498]) begin
            regVec_498 <= _zz_regVec_0;
          end
          if(_zz_1[499]) begin
            regVec_499 <= _zz_regVec_0;
          end
          if(_zz_1[500]) begin
            regVec_500 <= _zz_regVec_0;
          end
          if(_zz_1[501]) begin
            regVec_501 <= _zz_regVec_0;
          end
          if(_zz_1[502]) begin
            regVec_502 <= _zz_regVec_0;
          end
          if(_zz_1[503]) begin
            regVec_503 <= _zz_regVec_0;
          end
          if(_zz_1[504]) begin
            regVec_504 <= _zz_regVec_0;
          end
          if(_zz_1[505]) begin
            regVec_505 <= _zz_regVec_0;
          end
          if(_zz_1[506]) begin
            regVec_506 <= _zz_regVec_0;
          end
          if(_zz_1[507]) begin
            regVec_507 <= _zz_regVec_0;
          end
          if(_zz_1[508]) begin
            regVec_508 <= _zz_regVec_0;
          end
          if(_zz_1[509]) begin
            regVec_509 <= _zz_regVec_0;
          end
          if(_zz_1[510]) begin
            regVec_510 <= _zz_regVec_0;
          end
          if(_zz_1[511]) begin
            regVec_511 <= _zz_regVec_0;
          end
          if(_zz_1[512]) begin
            regVec_512 <= _zz_regVec_0;
          end
          if(_zz_1[513]) begin
            regVec_513 <= _zz_regVec_0;
          end
          if(_zz_1[514]) begin
            regVec_514 <= _zz_regVec_0;
          end
          if(_zz_1[515]) begin
            regVec_515 <= _zz_regVec_0;
          end
          if(_zz_1[516]) begin
            regVec_516 <= _zz_regVec_0;
          end
          if(_zz_1[517]) begin
            regVec_517 <= _zz_regVec_0;
          end
          if(_zz_1[518]) begin
            regVec_518 <= _zz_regVec_0;
          end
          if(_zz_1[519]) begin
            regVec_519 <= _zz_regVec_0;
          end
          if(_zz_1[520]) begin
            regVec_520 <= _zz_regVec_0;
          end
          if(_zz_1[521]) begin
            regVec_521 <= _zz_regVec_0;
          end
          if(_zz_1[522]) begin
            regVec_522 <= _zz_regVec_0;
          end
          if(_zz_1[523]) begin
            regVec_523 <= _zz_regVec_0;
          end
          if(_zz_1[524]) begin
            regVec_524 <= _zz_regVec_0;
          end
          if(_zz_1[525]) begin
            regVec_525 <= _zz_regVec_0;
          end
          if(_zz_1[526]) begin
            regVec_526 <= _zz_regVec_0;
          end
          if(_zz_1[527]) begin
            regVec_527 <= _zz_regVec_0;
          end
          if(_zz_1[528]) begin
            regVec_528 <= _zz_regVec_0;
          end
          if(_zz_1[529]) begin
            regVec_529 <= _zz_regVec_0;
          end
          if(_zz_1[530]) begin
            regVec_530 <= _zz_regVec_0;
          end
          if(_zz_1[531]) begin
            regVec_531 <= _zz_regVec_0;
          end
          if(_zz_1[532]) begin
            regVec_532 <= _zz_regVec_0;
          end
          if(_zz_1[533]) begin
            regVec_533 <= _zz_regVec_0;
          end
          if(_zz_1[534]) begin
            regVec_534 <= _zz_regVec_0;
          end
          if(_zz_1[535]) begin
            regVec_535 <= _zz_regVec_0;
          end
          if(_zz_1[536]) begin
            regVec_536 <= _zz_regVec_0;
          end
          if(_zz_1[537]) begin
            regVec_537 <= _zz_regVec_0;
          end
          if(_zz_1[538]) begin
            regVec_538 <= _zz_regVec_0;
          end
          if(_zz_1[539]) begin
            regVec_539 <= _zz_regVec_0;
          end
          if(_zz_1[540]) begin
            regVec_540 <= _zz_regVec_0;
          end
          if(_zz_1[541]) begin
            regVec_541 <= _zz_regVec_0;
          end
          if(_zz_1[542]) begin
            regVec_542 <= _zz_regVec_0;
          end
          if(_zz_1[543]) begin
            regVec_543 <= _zz_regVec_0;
          end
          if(_zz_1[544]) begin
            regVec_544 <= _zz_regVec_0;
          end
          if(_zz_1[545]) begin
            regVec_545 <= _zz_regVec_0;
          end
          if(_zz_1[546]) begin
            regVec_546 <= _zz_regVec_0;
          end
          if(_zz_1[547]) begin
            regVec_547 <= _zz_regVec_0;
          end
          if(_zz_1[548]) begin
            regVec_548 <= _zz_regVec_0;
          end
          if(_zz_1[549]) begin
            regVec_549 <= _zz_regVec_0;
          end
          if(_zz_1[550]) begin
            regVec_550 <= _zz_regVec_0;
          end
          if(_zz_1[551]) begin
            regVec_551 <= _zz_regVec_0;
          end
          if(_zz_1[552]) begin
            regVec_552 <= _zz_regVec_0;
          end
          if(_zz_1[553]) begin
            regVec_553 <= _zz_regVec_0;
          end
          if(_zz_1[554]) begin
            regVec_554 <= _zz_regVec_0;
          end
          if(_zz_1[555]) begin
            regVec_555 <= _zz_regVec_0;
          end
          if(_zz_1[556]) begin
            regVec_556 <= _zz_regVec_0;
          end
          if(_zz_1[557]) begin
            regVec_557 <= _zz_regVec_0;
          end
          if(_zz_1[558]) begin
            regVec_558 <= _zz_regVec_0;
          end
          if(_zz_1[559]) begin
            regVec_559 <= _zz_regVec_0;
          end
          if(_zz_1[560]) begin
            regVec_560 <= _zz_regVec_0;
          end
          if(_zz_1[561]) begin
            regVec_561 <= _zz_regVec_0;
          end
          if(_zz_1[562]) begin
            regVec_562 <= _zz_regVec_0;
          end
          if(_zz_1[563]) begin
            regVec_563 <= _zz_regVec_0;
          end
          if(_zz_1[564]) begin
            regVec_564 <= _zz_regVec_0;
          end
          if(_zz_1[565]) begin
            regVec_565 <= _zz_regVec_0;
          end
          if(_zz_1[566]) begin
            regVec_566 <= _zz_regVec_0;
          end
          if(_zz_1[567]) begin
            regVec_567 <= _zz_regVec_0;
          end
          if(_zz_1[568]) begin
            regVec_568 <= _zz_regVec_0;
          end
          if(_zz_1[569]) begin
            regVec_569 <= _zz_regVec_0;
          end
          if(_zz_1[570]) begin
            regVec_570 <= _zz_regVec_0;
          end
          if(_zz_1[571]) begin
            regVec_571 <= _zz_regVec_0;
          end
          if(_zz_1[572]) begin
            regVec_572 <= _zz_regVec_0;
          end
          if(_zz_1[573]) begin
            regVec_573 <= _zz_regVec_0;
          end
          if(_zz_1[574]) begin
            regVec_574 <= _zz_regVec_0;
          end
          if(_zz_1[575]) begin
            regVec_575 <= _zz_regVec_0;
          end
          if(_zz_1[576]) begin
            regVec_576 <= _zz_regVec_0;
          end
          if(_zz_1[577]) begin
            regVec_577 <= _zz_regVec_0;
          end
          if(_zz_1[578]) begin
            regVec_578 <= _zz_regVec_0;
          end
          if(_zz_1[579]) begin
            regVec_579 <= _zz_regVec_0;
          end
          if(_zz_1[580]) begin
            regVec_580 <= _zz_regVec_0;
          end
          if(_zz_1[581]) begin
            regVec_581 <= _zz_regVec_0;
          end
          if(_zz_1[582]) begin
            regVec_582 <= _zz_regVec_0;
          end
          if(_zz_1[583]) begin
            regVec_583 <= _zz_regVec_0;
          end
          if(_zz_1[584]) begin
            regVec_584 <= _zz_regVec_0;
          end
          if(_zz_1[585]) begin
            regVec_585 <= _zz_regVec_0;
          end
          if(_zz_1[586]) begin
            regVec_586 <= _zz_regVec_0;
          end
          if(_zz_1[587]) begin
            regVec_587 <= _zz_regVec_0;
          end
          if(_zz_1[588]) begin
            regVec_588 <= _zz_regVec_0;
          end
          if(_zz_1[589]) begin
            regVec_589 <= _zz_regVec_0;
          end
          if(_zz_1[590]) begin
            regVec_590 <= _zz_regVec_0;
          end
          if(_zz_1[591]) begin
            regVec_591 <= _zz_regVec_0;
          end
          if(_zz_1[592]) begin
            regVec_592 <= _zz_regVec_0;
          end
          if(_zz_1[593]) begin
            regVec_593 <= _zz_regVec_0;
          end
          if(_zz_1[594]) begin
            regVec_594 <= _zz_regVec_0;
          end
          if(_zz_1[595]) begin
            regVec_595 <= _zz_regVec_0;
          end
          if(_zz_1[596]) begin
            regVec_596 <= _zz_regVec_0;
          end
          if(_zz_1[597]) begin
            regVec_597 <= _zz_regVec_0;
          end
          if(_zz_1[598]) begin
            regVec_598 <= _zz_regVec_0;
          end
          if(_zz_1[599]) begin
            regVec_599 <= _zz_regVec_0;
          end
          if(_zz_1[600]) begin
            regVec_600 <= _zz_regVec_0;
          end
          if(_zz_1[601]) begin
            regVec_601 <= _zz_regVec_0;
          end
          if(_zz_1[602]) begin
            regVec_602 <= _zz_regVec_0;
          end
          if(_zz_1[603]) begin
            regVec_603 <= _zz_regVec_0;
          end
          if(_zz_1[604]) begin
            regVec_604 <= _zz_regVec_0;
          end
          if(_zz_1[605]) begin
            regVec_605 <= _zz_regVec_0;
          end
          if(_zz_1[606]) begin
            regVec_606 <= _zz_regVec_0;
          end
          if(_zz_1[607]) begin
            regVec_607 <= _zz_regVec_0;
          end
          if(_zz_1[608]) begin
            regVec_608 <= _zz_regVec_0;
          end
          if(_zz_1[609]) begin
            regVec_609 <= _zz_regVec_0;
          end
          if(_zz_1[610]) begin
            regVec_610 <= _zz_regVec_0;
          end
          if(_zz_1[611]) begin
            regVec_611 <= _zz_regVec_0;
          end
          if(_zz_1[612]) begin
            regVec_612 <= _zz_regVec_0;
          end
          if(_zz_1[613]) begin
            regVec_613 <= _zz_regVec_0;
          end
          if(_zz_1[614]) begin
            regVec_614 <= _zz_regVec_0;
          end
          if(_zz_1[615]) begin
            regVec_615 <= _zz_regVec_0;
          end
          if(_zz_1[616]) begin
            regVec_616 <= _zz_regVec_0;
          end
          if(_zz_1[617]) begin
            regVec_617 <= _zz_regVec_0;
          end
          if(_zz_1[618]) begin
            regVec_618 <= _zz_regVec_0;
          end
          if(_zz_1[619]) begin
            regVec_619 <= _zz_regVec_0;
          end
          if(_zz_1[620]) begin
            regVec_620 <= _zz_regVec_0;
          end
          if(_zz_1[621]) begin
            regVec_621 <= _zz_regVec_0;
          end
          if(_zz_1[622]) begin
            regVec_622 <= _zz_regVec_0;
          end
          if(_zz_1[623]) begin
            regVec_623 <= _zz_regVec_0;
          end
          if(_zz_1[624]) begin
            regVec_624 <= _zz_regVec_0;
          end
          if(_zz_1[625]) begin
            regVec_625 <= _zz_regVec_0;
          end
          if(_zz_1[626]) begin
            regVec_626 <= _zz_regVec_0;
          end
          if(_zz_1[627]) begin
            regVec_627 <= _zz_regVec_0;
          end
          if(_zz_1[628]) begin
            regVec_628 <= _zz_regVec_0;
          end
          if(_zz_1[629]) begin
            regVec_629 <= _zz_regVec_0;
          end
          if(_zz_1[630]) begin
            regVec_630 <= _zz_regVec_0;
          end
          if(_zz_1[631]) begin
            regVec_631 <= _zz_regVec_0;
          end
          if(_zz_1[632]) begin
            regVec_632 <= _zz_regVec_0;
          end
          if(_zz_1[633]) begin
            regVec_633 <= _zz_regVec_0;
          end
          if(_zz_1[634]) begin
            regVec_634 <= _zz_regVec_0;
          end
          if(_zz_1[635]) begin
            regVec_635 <= _zz_regVec_0;
          end
          if(_zz_1[636]) begin
            regVec_636 <= _zz_regVec_0;
          end
          if(_zz_1[637]) begin
            regVec_637 <= _zz_regVec_0;
          end
          if(_zz_1[638]) begin
            regVec_638 <= _zz_regVec_0;
          end
          if(_zz_1[639]) begin
            regVec_639 <= _zz_regVec_0;
          end
          if(_zz_1[640]) begin
            regVec_640 <= _zz_regVec_0;
          end
          if(_zz_1[641]) begin
            regVec_641 <= _zz_regVec_0;
          end
          if(_zz_1[642]) begin
            regVec_642 <= _zz_regVec_0;
          end
          if(_zz_1[643]) begin
            regVec_643 <= _zz_regVec_0;
          end
          if(_zz_1[644]) begin
            regVec_644 <= _zz_regVec_0;
          end
          if(_zz_1[645]) begin
            regVec_645 <= _zz_regVec_0;
          end
          if(_zz_1[646]) begin
            regVec_646 <= _zz_regVec_0;
          end
          if(_zz_1[647]) begin
            regVec_647 <= _zz_regVec_0;
          end
          if(_zz_1[648]) begin
            regVec_648 <= _zz_regVec_0;
          end
          if(_zz_1[649]) begin
            regVec_649 <= _zz_regVec_0;
          end
          if(_zz_1[650]) begin
            regVec_650 <= _zz_regVec_0;
          end
          if(_zz_1[651]) begin
            regVec_651 <= _zz_regVec_0;
          end
          if(_zz_1[652]) begin
            regVec_652 <= _zz_regVec_0;
          end
          if(_zz_1[653]) begin
            regVec_653 <= _zz_regVec_0;
          end
          if(_zz_1[654]) begin
            regVec_654 <= _zz_regVec_0;
          end
          if(_zz_1[655]) begin
            regVec_655 <= _zz_regVec_0;
          end
          if(_zz_1[656]) begin
            regVec_656 <= _zz_regVec_0;
          end
          if(_zz_1[657]) begin
            regVec_657 <= _zz_regVec_0;
          end
          if(_zz_1[658]) begin
            regVec_658 <= _zz_regVec_0;
          end
          if(_zz_1[659]) begin
            regVec_659 <= _zz_regVec_0;
          end
          if(_zz_1[660]) begin
            regVec_660 <= _zz_regVec_0;
          end
          if(_zz_1[661]) begin
            regVec_661 <= _zz_regVec_0;
          end
          if(_zz_1[662]) begin
            regVec_662 <= _zz_regVec_0;
          end
          if(_zz_1[663]) begin
            regVec_663 <= _zz_regVec_0;
          end
          if(_zz_1[664]) begin
            regVec_664 <= _zz_regVec_0;
          end
          if(_zz_1[665]) begin
            regVec_665 <= _zz_regVec_0;
          end
          if(_zz_1[666]) begin
            regVec_666 <= _zz_regVec_0;
          end
          if(_zz_1[667]) begin
            regVec_667 <= _zz_regVec_0;
          end
          if(_zz_1[668]) begin
            regVec_668 <= _zz_regVec_0;
          end
          if(_zz_1[669]) begin
            regVec_669 <= _zz_regVec_0;
          end
          if(_zz_1[670]) begin
            regVec_670 <= _zz_regVec_0;
          end
          if(_zz_1[671]) begin
            regVec_671 <= _zz_regVec_0;
          end
          if(_zz_1[672]) begin
            regVec_672 <= _zz_regVec_0;
          end
          if(_zz_1[673]) begin
            regVec_673 <= _zz_regVec_0;
          end
          if(_zz_1[674]) begin
            regVec_674 <= _zz_regVec_0;
          end
          if(_zz_1[675]) begin
            regVec_675 <= _zz_regVec_0;
          end
          if(_zz_1[676]) begin
            regVec_676 <= _zz_regVec_0;
          end
          if(_zz_1[677]) begin
            regVec_677 <= _zz_regVec_0;
          end
          if(_zz_1[678]) begin
            regVec_678 <= _zz_regVec_0;
          end
          if(_zz_1[679]) begin
            regVec_679 <= _zz_regVec_0;
          end
          if(_zz_1[680]) begin
            regVec_680 <= _zz_regVec_0;
          end
          if(_zz_1[681]) begin
            regVec_681 <= _zz_regVec_0;
          end
          if(_zz_1[682]) begin
            regVec_682 <= _zz_regVec_0;
          end
          if(_zz_1[683]) begin
            regVec_683 <= _zz_regVec_0;
          end
          if(_zz_1[684]) begin
            regVec_684 <= _zz_regVec_0;
          end
          if(_zz_1[685]) begin
            regVec_685 <= _zz_regVec_0;
          end
          if(_zz_1[686]) begin
            regVec_686 <= _zz_regVec_0;
          end
          if(_zz_1[687]) begin
            regVec_687 <= _zz_regVec_0;
          end
          if(_zz_1[688]) begin
            regVec_688 <= _zz_regVec_0;
          end
          if(_zz_1[689]) begin
            regVec_689 <= _zz_regVec_0;
          end
          if(_zz_1[690]) begin
            regVec_690 <= _zz_regVec_0;
          end
          if(_zz_1[691]) begin
            regVec_691 <= _zz_regVec_0;
          end
          if(_zz_1[692]) begin
            regVec_692 <= _zz_regVec_0;
          end
          if(_zz_1[693]) begin
            regVec_693 <= _zz_regVec_0;
          end
          if(_zz_1[694]) begin
            regVec_694 <= _zz_regVec_0;
          end
          if(_zz_1[695]) begin
            regVec_695 <= _zz_regVec_0;
          end
          if(_zz_1[696]) begin
            regVec_696 <= _zz_regVec_0;
          end
          if(_zz_1[697]) begin
            regVec_697 <= _zz_regVec_0;
          end
          if(_zz_1[698]) begin
            regVec_698 <= _zz_regVec_0;
          end
          if(_zz_1[699]) begin
            regVec_699 <= _zz_regVec_0;
          end
          if(_zz_1[700]) begin
            regVec_700 <= _zz_regVec_0;
          end
          if(_zz_1[701]) begin
            regVec_701 <= _zz_regVec_0;
          end
          if(_zz_1[702]) begin
            regVec_702 <= _zz_regVec_0;
          end
          if(_zz_1[703]) begin
            regVec_703 <= _zz_regVec_0;
          end
          if(_zz_1[704]) begin
            regVec_704 <= _zz_regVec_0;
          end
          if(_zz_1[705]) begin
            regVec_705 <= _zz_regVec_0;
          end
          if(_zz_1[706]) begin
            regVec_706 <= _zz_regVec_0;
          end
          if(_zz_1[707]) begin
            regVec_707 <= _zz_regVec_0;
          end
          if(_zz_1[708]) begin
            regVec_708 <= _zz_regVec_0;
          end
          if(_zz_1[709]) begin
            regVec_709 <= _zz_regVec_0;
          end
          if(_zz_1[710]) begin
            regVec_710 <= _zz_regVec_0;
          end
          if(_zz_1[711]) begin
            regVec_711 <= _zz_regVec_0;
          end
          if(_zz_1[712]) begin
            regVec_712 <= _zz_regVec_0;
          end
          if(_zz_1[713]) begin
            regVec_713 <= _zz_regVec_0;
          end
          if(_zz_1[714]) begin
            regVec_714 <= _zz_regVec_0;
          end
          if(_zz_1[715]) begin
            regVec_715 <= _zz_regVec_0;
          end
          if(_zz_1[716]) begin
            regVec_716 <= _zz_regVec_0;
          end
          if(_zz_1[717]) begin
            regVec_717 <= _zz_regVec_0;
          end
          if(_zz_1[718]) begin
            regVec_718 <= _zz_regVec_0;
          end
          if(_zz_1[719]) begin
            regVec_719 <= _zz_regVec_0;
          end
          if(_zz_1[720]) begin
            regVec_720 <= _zz_regVec_0;
          end
          if(_zz_1[721]) begin
            regVec_721 <= _zz_regVec_0;
          end
          if(_zz_1[722]) begin
            regVec_722 <= _zz_regVec_0;
          end
          if(_zz_1[723]) begin
            regVec_723 <= _zz_regVec_0;
          end
          if(_zz_1[724]) begin
            regVec_724 <= _zz_regVec_0;
          end
          if(_zz_1[725]) begin
            regVec_725 <= _zz_regVec_0;
          end
          if(_zz_1[726]) begin
            regVec_726 <= _zz_regVec_0;
          end
          if(_zz_1[727]) begin
            regVec_727 <= _zz_regVec_0;
          end
          if(_zz_1[728]) begin
            regVec_728 <= _zz_regVec_0;
          end
          if(_zz_1[729]) begin
            regVec_729 <= _zz_regVec_0;
          end
          if(_zz_1[730]) begin
            regVec_730 <= _zz_regVec_0;
          end
          if(_zz_1[731]) begin
            regVec_731 <= _zz_regVec_0;
          end
          if(_zz_1[732]) begin
            regVec_732 <= _zz_regVec_0;
          end
          if(_zz_1[733]) begin
            regVec_733 <= _zz_regVec_0;
          end
          if(_zz_1[734]) begin
            regVec_734 <= _zz_regVec_0;
          end
          if(_zz_1[735]) begin
            regVec_735 <= _zz_regVec_0;
          end
          if(_zz_1[736]) begin
            regVec_736 <= _zz_regVec_0;
          end
          if(_zz_1[737]) begin
            regVec_737 <= _zz_regVec_0;
          end
          if(_zz_1[738]) begin
            regVec_738 <= _zz_regVec_0;
          end
          if(_zz_1[739]) begin
            regVec_739 <= _zz_regVec_0;
          end
          if(_zz_1[740]) begin
            regVec_740 <= _zz_regVec_0;
          end
          if(_zz_1[741]) begin
            regVec_741 <= _zz_regVec_0;
          end
          if(_zz_1[742]) begin
            regVec_742 <= _zz_regVec_0;
          end
          if(_zz_1[743]) begin
            regVec_743 <= _zz_regVec_0;
          end
          if(_zz_1[744]) begin
            regVec_744 <= _zz_regVec_0;
          end
          if(_zz_1[745]) begin
            regVec_745 <= _zz_regVec_0;
          end
          if(_zz_1[746]) begin
            regVec_746 <= _zz_regVec_0;
          end
          if(_zz_1[747]) begin
            regVec_747 <= _zz_regVec_0;
          end
          if(_zz_1[748]) begin
            regVec_748 <= _zz_regVec_0;
          end
          if(_zz_1[749]) begin
            regVec_749 <= _zz_regVec_0;
          end
          if(_zz_1[750]) begin
            regVec_750 <= _zz_regVec_0;
          end
          if(_zz_1[751]) begin
            regVec_751 <= _zz_regVec_0;
          end
          if(_zz_1[752]) begin
            regVec_752 <= _zz_regVec_0;
          end
          if(_zz_1[753]) begin
            regVec_753 <= _zz_regVec_0;
          end
          if(_zz_1[754]) begin
            regVec_754 <= _zz_regVec_0;
          end
          if(_zz_1[755]) begin
            regVec_755 <= _zz_regVec_0;
          end
          if(_zz_1[756]) begin
            regVec_756 <= _zz_regVec_0;
          end
          if(_zz_1[757]) begin
            regVec_757 <= _zz_regVec_0;
          end
          if(_zz_1[758]) begin
            regVec_758 <= _zz_regVec_0;
          end
          if(_zz_1[759]) begin
            regVec_759 <= _zz_regVec_0;
          end
          if(_zz_1[760]) begin
            regVec_760 <= _zz_regVec_0;
          end
          if(_zz_1[761]) begin
            regVec_761 <= _zz_regVec_0;
          end
          if(_zz_1[762]) begin
            regVec_762 <= _zz_regVec_0;
          end
          if(_zz_1[763]) begin
            regVec_763 <= _zz_regVec_0;
          end
          if(_zz_1[764]) begin
            regVec_764 <= _zz_regVec_0;
          end
          if(_zz_1[765]) begin
            regVec_765 <= _zz_regVec_0;
          end
          if(_zz_1[766]) begin
            regVec_766 <= _zz_regVec_0;
          end
          if(_zz_1[767]) begin
            regVec_767 <= _zz_regVec_0;
          end
          if(_zz_1[768]) begin
            regVec_768 <= _zz_regVec_0;
          end
          if(_zz_1[769]) begin
            regVec_769 <= _zz_regVec_0;
          end
          if(_zz_1[770]) begin
            regVec_770 <= _zz_regVec_0;
          end
          if(_zz_1[771]) begin
            regVec_771 <= _zz_regVec_0;
          end
          if(_zz_1[772]) begin
            regVec_772 <= _zz_regVec_0;
          end
          if(_zz_1[773]) begin
            regVec_773 <= _zz_regVec_0;
          end
          if(_zz_1[774]) begin
            regVec_774 <= _zz_regVec_0;
          end
          if(_zz_1[775]) begin
            regVec_775 <= _zz_regVec_0;
          end
          if(_zz_1[776]) begin
            regVec_776 <= _zz_regVec_0;
          end
          if(_zz_1[777]) begin
            regVec_777 <= _zz_regVec_0;
          end
          if(_zz_1[778]) begin
            regVec_778 <= _zz_regVec_0;
          end
          if(_zz_1[779]) begin
            regVec_779 <= _zz_regVec_0;
          end
          if(_zz_1[780]) begin
            regVec_780 <= _zz_regVec_0;
          end
          if(_zz_1[781]) begin
            regVec_781 <= _zz_regVec_0;
          end
          if(_zz_1[782]) begin
            regVec_782 <= _zz_regVec_0;
          end
          if(_zz_1[783]) begin
            regVec_783 <= _zz_regVec_0;
          end
          if(_zz_1[784]) begin
            regVec_784 <= _zz_regVec_0;
          end
          if(_zz_1[785]) begin
            regVec_785 <= _zz_regVec_0;
          end
          if(_zz_1[786]) begin
            regVec_786 <= _zz_regVec_0;
          end
          if(_zz_1[787]) begin
            regVec_787 <= _zz_regVec_0;
          end
          if(_zz_1[788]) begin
            regVec_788 <= _zz_regVec_0;
          end
          if(_zz_1[789]) begin
            regVec_789 <= _zz_regVec_0;
          end
          if(_zz_1[790]) begin
            regVec_790 <= _zz_regVec_0;
          end
          if(_zz_1[791]) begin
            regVec_791 <= _zz_regVec_0;
          end
          if(_zz_1[792]) begin
            regVec_792 <= _zz_regVec_0;
          end
          if(_zz_1[793]) begin
            regVec_793 <= _zz_regVec_0;
          end
          if(_zz_1[794]) begin
            regVec_794 <= _zz_regVec_0;
          end
          if(_zz_1[795]) begin
            regVec_795 <= _zz_regVec_0;
          end
          if(_zz_1[796]) begin
            regVec_796 <= _zz_regVec_0;
          end
          if(_zz_1[797]) begin
            regVec_797 <= _zz_regVec_0;
          end
          if(_zz_1[798]) begin
            regVec_798 <= _zz_regVec_0;
          end
          if(_zz_1[799]) begin
            regVec_799 <= _zz_regVec_0;
          end
          if(_zz_1[800]) begin
            regVec_800 <= _zz_regVec_0;
          end
          if(_zz_1[801]) begin
            regVec_801 <= _zz_regVec_0;
          end
          if(_zz_1[802]) begin
            regVec_802 <= _zz_regVec_0;
          end
          if(_zz_1[803]) begin
            regVec_803 <= _zz_regVec_0;
          end
          if(_zz_1[804]) begin
            regVec_804 <= _zz_regVec_0;
          end
          if(_zz_1[805]) begin
            regVec_805 <= _zz_regVec_0;
          end
          if(_zz_1[806]) begin
            regVec_806 <= _zz_regVec_0;
          end
          if(_zz_1[807]) begin
            regVec_807 <= _zz_regVec_0;
          end
          if(_zz_1[808]) begin
            regVec_808 <= _zz_regVec_0;
          end
          if(_zz_1[809]) begin
            regVec_809 <= _zz_regVec_0;
          end
          if(_zz_1[810]) begin
            regVec_810 <= _zz_regVec_0;
          end
          if(_zz_1[811]) begin
            regVec_811 <= _zz_regVec_0;
          end
          if(_zz_1[812]) begin
            regVec_812 <= _zz_regVec_0;
          end
          if(_zz_1[813]) begin
            regVec_813 <= _zz_regVec_0;
          end
          if(_zz_1[814]) begin
            regVec_814 <= _zz_regVec_0;
          end
          if(_zz_1[815]) begin
            regVec_815 <= _zz_regVec_0;
          end
          if(_zz_1[816]) begin
            regVec_816 <= _zz_regVec_0;
          end
          if(_zz_1[817]) begin
            regVec_817 <= _zz_regVec_0;
          end
          if(_zz_1[818]) begin
            regVec_818 <= _zz_regVec_0;
          end
          if(_zz_1[819]) begin
            regVec_819 <= _zz_regVec_0;
          end
          if(_zz_1[820]) begin
            regVec_820 <= _zz_regVec_0;
          end
          if(_zz_1[821]) begin
            regVec_821 <= _zz_regVec_0;
          end
          if(_zz_1[822]) begin
            regVec_822 <= _zz_regVec_0;
          end
          if(_zz_1[823]) begin
            regVec_823 <= _zz_regVec_0;
          end
          if(_zz_1[824]) begin
            regVec_824 <= _zz_regVec_0;
          end
          if(_zz_1[825]) begin
            regVec_825 <= _zz_regVec_0;
          end
          if(_zz_1[826]) begin
            regVec_826 <= _zz_regVec_0;
          end
          if(_zz_1[827]) begin
            regVec_827 <= _zz_regVec_0;
          end
          if(_zz_1[828]) begin
            regVec_828 <= _zz_regVec_0;
          end
          if(_zz_1[829]) begin
            regVec_829 <= _zz_regVec_0;
          end
          if(_zz_1[830]) begin
            regVec_830 <= _zz_regVec_0;
          end
          if(_zz_1[831]) begin
            regVec_831 <= _zz_regVec_0;
          end
          if(_zz_1[832]) begin
            regVec_832 <= _zz_regVec_0;
          end
          if(_zz_1[833]) begin
            regVec_833 <= _zz_regVec_0;
          end
          if(_zz_1[834]) begin
            regVec_834 <= _zz_regVec_0;
          end
          if(_zz_1[835]) begin
            regVec_835 <= _zz_regVec_0;
          end
          if(_zz_1[836]) begin
            regVec_836 <= _zz_regVec_0;
          end
          if(_zz_1[837]) begin
            regVec_837 <= _zz_regVec_0;
          end
          if(_zz_1[838]) begin
            regVec_838 <= _zz_regVec_0;
          end
          if(_zz_1[839]) begin
            regVec_839 <= _zz_regVec_0;
          end
          if(_zz_1[840]) begin
            regVec_840 <= _zz_regVec_0;
          end
          if(_zz_1[841]) begin
            regVec_841 <= _zz_regVec_0;
          end
          if(_zz_1[842]) begin
            regVec_842 <= _zz_regVec_0;
          end
          if(_zz_1[843]) begin
            regVec_843 <= _zz_regVec_0;
          end
          if(_zz_1[844]) begin
            regVec_844 <= _zz_regVec_0;
          end
          if(_zz_1[845]) begin
            regVec_845 <= _zz_regVec_0;
          end
          if(_zz_1[846]) begin
            regVec_846 <= _zz_regVec_0;
          end
          if(_zz_1[847]) begin
            regVec_847 <= _zz_regVec_0;
          end
          if(_zz_1[848]) begin
            regVec_848 <= _zz_regVec_0;
          end
          if(_zz_1[849]) begin
            regVec_849 <= _zz_regVec_0;
          end
          if(_zz_1[850]) begin
            regVec_850 <= _zz_regVec_0;
          end
          if(_zz_1[851]) begin
            regVec_851 <= _zz_regVec_0;
          end
          if(_zz_1[852]) begin
            regVec_852 <= _zz_regVec_0;
          end
          if(_zz_1[853]) begin
            regVec_853 <= _zz_regVec_0;
          end
          if(_zz_1[854]) begin
            regVec_854 <= _zz_regVec_0;
          end
          if(_zz_1[855]) begin
            regVec_855 <= _zz_regVec_0;
          end
          if(_zz_1[856]) begin
            regVec_856 <= _zz_regVec_0;
          end
          if(_zz_1[857]) begin
            regVec_857 <= _zz_regVec_0;
          end
          if(_zz_1[858]) begin
            regVec_858 <= _zz_regVec_0;
          end
          if(_zz_1[859]) begin
            regVec_859 <= _zz_regVec_0;
          end
          if(_zz_1[860]) begin
            regVec_860 <= _zz_regVec_0;
          end
          if(_zz_1[861]) begin
            regVec_861 <= _zz_regVec_0;
          end
          if(_zz_1[862]) begin
            regVec_862 <= _zz_regVec_0;
          end
          if(_zz_1[863]) begin
            regVec_863 <= _zz_regVec_0;
          end
          if(_zz_1[864]) begin
            regVec_864 <= _zz_regVec_0;
          end
          if(_zz_1[865]) begin
            regVec_865 <= _zz_regVec_0;
          end
          if(_zz_1[866]) begin
            regVec_866 <= _zz_regVec_0;
          end
          if(_zz_1[867]) begin
            regVec_867 <= _zz_regVec_0;
          end
          if(_zz_1[868]) begin
            regVec_868 <= _zz_regVec_0;
          end
          if(_zz_1[869]) begin
            regVec_869 <= _zz_regVec_0;
          end
          if(_zz_1[870]) begin
            regVec_870 <= _zz_regVec_0;
          end
          if(_zz_1[871]) begin
            regVec_871 <= _zz_regVec_0;
          end
          if(_zz_1[872]) begin
            regVec_872 <= _zz_regVec_0;
          end
          if(_zz_1[873]) begin
            regVec_873 <= _zz_regVec_0;
          end
          if(_zz_1[874]) begin
            regVec_874 <= _zz_regVec_0;
          end
          if(_zz_1[875]) begin
            regVec_875 <= _zz_regVec_0;
          end
          if(_zz_1[876]) begin
            regVec_876 <= _zz_regVec_0;
          end
          if(_zz_1[877]) begin
            regVec_877 <= _zz_regVec_0;
          end
          if(_zz_1[878]) begin
            regVec_878 <= _zz_regVec_0;
          end
          if(_zz_1[879]) begin
            regVec_879 <= _zz_regVec_0;
          end
          if(_zz_1[880]) begin
            regVec_880 <= _zz_regVec_0;
          end
          if(_zz_1[881]) begin
            regVec_881 <= _zz_regVec_0;
          end
          if(_zz_1[882]) begin
            regVec_882 <= _zz_regVec_0;
          end
          if(_zz_1[883]) begin
            regVec_883 <= _zz_regVec_0;
          end
          if(_zz_1[884]) begin
            regVec_884 <= _zz_regVec_0;
          end
          if(_zz_1[885]) begin
            regVec_885 <= _zz_regVec_0;
          end
          if(_zz_1[886]) begin
            regVec_886 <= _zz_regVec_0;
          end
          if(_zz_1[887]) begin
            regVec_887 <= _zz_regVec_0;
          end
          if(_zz_1[888]) begin
            regVec_888 <= _zz_regVec_0;
          end
          if(_zz_1[889]) begin
            regVec_889 <= _zz_regVec_0;
          end
          if(_zz_1[890]) begin
            regVec_890 <= _zz_regVec_0;
          end
          if(_zz_1[891]) begin
            regVec_891 <= _zz_regVec_0;
          end
          if(_zz_1[892]) begin
            regVec_892 <= _zz_regVec_0;
          end
          if(_zz_1[893]) begin
            regVec_893 <= _zz_regVec_0;
          end
          if(_zz_1[894]) begin
            regVec_894 <= _zz_regVec_0;
          end
          if(_zz_1[895]) begin
            regVec_895 <= _zz_regVec_0;
          end
          if(_zz_1[896]) begin
            regVec_896 <= _zz_regVec_0;
          end
          if(_zz_1[897]) begin
            regVec_897 <= _zz_regVec_0;
          end
          if(_zz_1[898]) begin
            regVec_898 <= _zz_regVec_0;
          end
          if(_zz_1[899]) begin
            regVec_899 <= _zz_regVec_0;
          end
          if(_zz_1[900]) begin
            regVec_900 <= _zz_regVec_0;
          end
          if(_zz_1[901]) begin
            regVec_901 <= _zz_regVec_0;
          end
          if(_zz_1[902]) begin
            regVec_902 <= _zz_regVec_0;
          end
          if(_zz_1[903]) begin
            regVec_903 <= _zz_regVec_0;
          end
          if(_zz_1[904]) begin
            regVec_904 <= _zz_regVec_0;
          end
          if(_zz_1[905]) begin
            regVec_905 <= _zz_regVec_0;
          end
          if(_zz_1[906]) begin
            regVec_906 <= _zz_regVec_0;
          end
          if(_zz_1[907]) begin
            regVec_907 <= _zz_regVec_0;
          end
          if(_zz_1[908]) begin
            regVec_908 <= _zz_regVec_0;
          end
          if(_zz_1[909]) begin
            regVec_909 <= _zz_regVec_0;
          end
          if(_zz_1[910]) begin
            regVec_910 <= _zz_regVec_0;
          end
          if(_zz_1[911]) begin
            regVec_911 <= _zz_regVec_0;
          end
          if(_zz_1[912]) begin
            regVec_912 <= _zz_regVec_0;
          end
          if(_zz_1[913]) begin
            regVec_913 <= _zz_regVec_0;
          end
          if(_zz_1[914]) begin
            regVec_914 <= _zz_regVec_0;
          end
          if(_zz_1[915]) begin
            regVec_915 <= _zz_regVec_0;
          end
          if(_zz_1[916]) begin
            regVec_916 <= _zz_regVec_0;
          end
          if(_zz_1[917]) begin
            regVec_917 <= _zz_regVec_0;
          end
          if(_zz_1[918]) begin
            regVec_918 <= _zz_regVec_0;
          end
          if(_zz_1[919]) begin
            regVec_919 <= _zz_regVec_0;
          end
          if(_zz_1[920]) begin
            regVec_920 <= _zz_regVec_0;
          end
          if(_zz_1[921]) begin
            regVec_921 <= _zz_regVec_0;
          end
          if(_zz_1[922]) begin
            regVec_922 <= _zz_regVec_0;
          end
          if(_zz_1[923]) begin
            regVec_923 <= _zz_regVec_0;
          end
          if(_zz_1[924]) begin
            regVec_924 <= _zz_regVec_0;
          end
          if(_zz_1[925]) begin
            regVec_925 <= _zz_regVec_0;
          end
          if(_zz_1[926]) begin
            regVec_926 <= _zz_regVec_0;
          end
          if(_zz_1[927]) begin
            regVec_927 <= _zz_regVec_0;
          end
          if(_zz_1[928]) begin
            regVec_928 <= _zz_regVec_0;
          end
          if(_zz_1[929]) begin
            regVec_929 <= _zz_regVec_0;
          end
          if(_zz_1[930]) begin
            regVec_930 <= _zz_regVec_0;
          end
          if(_zz_1[931]) begin
            regVec_931 <= _zz_regVec_0;
          end
          if(_zz_1[932]) begin
            regVec_932 <= _zz_regVec_0;
          end
          if(_zz_1[933]) begin
            regVec_933 <= _zz_regVec_0;
          end
          if(_zz_1[934]) begin
            regVec_934 <= _zz_regVec_0;
          end
          if(_zz_1[935]) begin
            regVec_935 <= _zz_regVec_0;
          end
          if(_zz_1[936]) begin
            regVec_936 <= _zz_regVec_0;
          end
          if(_zz_1[937]) begin
            regVec_937 <= _zz_regVec_0;
          end
          if(_zz_1[938]) begin
            regVec_938 <= _zz_regVec_0;
          end
          if(_zz_1[939]) begin
            regVec_939 <= _zz_regVec_0;
          end
          if(_zz_1[940]) begin
            regVec_940 <= _zz_regVec_0;
          end
          if(_zz_1[941]) begin
            regVec_941 <= _zz_regVec_0;
          end
          if(_zz_1[942]) begin
            regVec_942 <= _zz_regVec_0;
          end
          if(_zz_1[943]) begin
            regVec_943 <= _zz_regVec_0;
          end
          if(_zz_1[944]) begin
            regVec_944 <= _zz_regVec_0;
          end
          if(_zz_1[945]) begin
            regVec_945 <= _zz_regVec_0;
          end
          if(_zz_1[946]) begin
            regVec_946 <= _zz_regVec_0;
          end
          if(_zz_1[947]) begin
            regVec_947 <= _zz_regVec_0;
          end
          if(_zz_1[948]) begin
            regVec_948 <= _zz_regVec_0;
          end
          if(_zz_1[949]) begin
            regVec_949 <= _zz_regVec_0;
          end
          if(_zz_1[950]) begin
            regVec_950 <= _zz_regVec_0;
          end
          if(_zz_1[951]) begin
            regVec_951 <= _zz_regVec_0;
          end
          if(_zz_1[952]) begin
            regVec_952 <= _zz_regVec_0;
          end
          if(_zz_1[953]) begin
            regVec_953 <= _zz_regVec_0;
          end
          if(_zz_1[954]) begin
            regVec_954 <= _zz_regVec_0;
          end
          if(_zz_1[955]) begin
            regVec_955 <= _zz_regVec_0;
          end
          if(_zz_1[956]) begin
            regVec_956 <= _zz_regVec_0;
          end
          if(_zz_1[957]) begin
            regVec_957 <= _zz_regVec_0;
          end
          if(_zz_1[958]) begin
            regVec_958 <= _zz_regVec_0;
          end
          if(_zz_1[959]) begin
            regVec_959 <= _zz_regVec_0;
          end
          if(_zz_1[960]) begin
            regVec_960 <= _zz_regVec_0;
          end
          if(_zz_1[961]) begin
            regVec_961 <= _zz_regVec_0;
          end
          if(_zz_1[962]) begin
            regVec_962 <= _zz_regVec_0;
          end
          if(_zz_1[963]) begin
            regVec_963 <= _zz_regVec_0;
          end
          if(_zz_1[964]) begin
            regVec_964 <= _zz_regVec_0;
          end
          if(_zz_1[965]) begin
            regVec_965 <= _zz_regVec_0;
          end
          if(_zz_1[966]) begin
            regVec_966 <= _zz_regVec_0;
          end
          if(_zz_1[967]) begin
            regVec_967 <= _zz_regVec_0;
          end
          if(_zz_1[968]) begin
            regVec_968 <= _zz_regVec_0;
          end
          if(_zz_1[969]) begin
            regVec_969 <= _zz_regVec_0;
          end
          if(_zz_1[970]) begin
            regVec_970 <= _zz_regVec_0;
          end
          if(_zz_1[971]) begin
            regVec_971 <= _zz_regVec_0;
          end
          if(_zz_1[972]) begin
            regVec_972 <= _zz_regVec_0;
          end
          if(_zz_1[973]) begin
            regVec_973 <= _zz_regVec_0;
          end
          if(_zz_1[974]) begin
            regVec_974 <= _zz_regVec_0;
          end
          if(_zz_1[975]) begin
            regVec_975 <= _zz_regVec_0;
          end
          if(_zz_1[976]) begin
            regVec_976 <= _zz_regVec_0;
          end
          if(_zz_1[977]) begin
            regVec_977 <= _zz_regVec_0;
          end
          if(_zz_1[978]) begin
            regVec_978 <= _zz_regVec_0;
          end
          if(_zz_1[979]) begin
            regVec_979 <= _zz_regVec_0;
          end
          if(_zz_1[980]) begin
            regVec_980 <= _zz_regVec_0;
          end
          if(_zz_1[981]) begin
            regVec_981 <= _zz_regVec_0;
          end
          if(_zz_1[982]) begin
            regVec_982 <= _zz_regVec_0;
          end
          if(_zz_1[983]) begin
            regVec_983 <= _zz_regVec_0;
          end
          if(_zz_1[984]) begin
            regVec_984 <= _zz_regVec_0;
          end
          if(_zz_1[985]) begin
            regVec_985 <= _zz_regVec_0;
          end
          if(_zz_1[986]) begin
            regVec_986 <= _zz_regVec_0;
          end
          if(_zz_1[987]) begin
            regVec_987 <= _zz_regVec_0;
          end
          if(_zz_1[988]) begin
            regVec_988 <= _zz_regVec_0;
          end
          if(_zz_1[989]) begin
            regVec_989 <= _zz_regVec_0;
          end
          if(_zz_1[990]) begin
            regVec_990 <= _zz_regVec_0;
          end
          if(_zz_1[991]) begin
            regVec_991 <= _zz_regVec_0;
          end
          if(_zz_1[992]) begin
            regVec_992 <= _zz_regVec_0;
          end
          if(_zz_1[993]) begin
            regVec_993 <= _zz_regVec_0;
          end
          if(_zz_1[994]) begin
            regVec_994 <= _zz_regVec_0;
          end
          if(_zz_1[995]) begin
            regVec_995 <= _zz_regVec_0;
          end
          if(_zz_1[996]) begin
            regVec_996 <= _zz_regVec_0;
          end
          if(_zz_1[997]) begin
            regVec_997 <= _zz_regVec_0;
          end
          if(_zz_1[998]) begin
            regVec_998 <= _zz_regVec_0;
          end
          if(_zz_1[999]) begin
            regVec_999 <= _zz_regVec_0;
          end
          if(_zz_1[1000]) begin
            regVec_1000 <= _zz_regVec_0;
          end
          if(_zz_1[1001]) begin
            regVec_1001 <= _zz_regVec_0;
          end
          if(_zz_1[1002]) begin
            regVec_1002 <= _zz_regVec_0;
          end
          if(_zz_1[1003]) begin
            regVec_1003 <= _zz_regVec_0;
          end
          if(_zz_1[1004]) begin
            regVec_1004 <= _zz_regVec_0;
          end
          if(_zz_1[1005]) begin
            regVec_1005 <= _zz_regVec_0;
          end
          if(_zz_1[1006]) begin
            regVec_1006 <= _zz_regVec_0;
          end
          if(_zz_1[1007]) begin
            regVec_1007 <= _zz_regVec_0;
          end
          if(_zz_1[1008]) begin
            regVec_1008 <= _zz_regVec_0;
          end
          if(_zz_1[1009]) begin
            regVec_1009 <= _zz_regVec_0;
          end
          if(_zz_1[1010]) begin
            regVec_1010 <= _zz_regVec_0;
          end
          if(_zz_1[1011]) begin
            regVec_1011 <= _zz_regVec_0;
          end
          if(_zz_1[1012]) begin
            regVec_1012 <= _zz_regVec_0;
          end
          if(_zz_1[1013]) begin
            regVec_1013 <= _zz_regVec_0;
          end
          if(_zz_1[1014]) begin
            regVec_1014 <= _zz_regVec_0;
          end
          if(_zz_1[1015]) begin
            regVec_1015 <= _zz_regVec_0;
          end
          if(_zz_1[1016]) begin
            regVec_1016 <= _zz_regVec_0;
          end
          if(_zz_1[1017]) begin
            regVec_1017 <= _zz_regVec_0;
          end
          if(_zz_1[1018]) begin
            regVec_1018 <= _zz_regVec_0;
          end
          if(_zz_1[1019]) begin
            regVec_1019 <= _zz_regVec_0;
          end
          if(_zz_1[1020]) begin
            regVec_1020 <= _zz_regVec_0;
          end
          if(_zz_1[1021]) begin
            regVec_1021 <= _zz_regVec_0;
          end
          if(_zz_1[1022]) begin
            regVec_1022 <= _zz_regVec_0;
          end
          if(_zz_1[1023]) begin
            regVec_1023 <= _zz_regVec_0;
          end
          if(_zz_1[1024]) begin
            regVec_1024 <= _zz_regVec_0;
          end
          if(_zz_1[1025]) begin
            regVec_1025 <= _zz_regVec_0;
          end
          if(_zz_1[1026]) begin
            regVec_1026 <= _zz_regVec_0;
          end
          if(_zz_1[1027]) begin
            regVec_1027 <= _zz_regVec_0;
          end
          if(_zz_1[1028]) begin
            regVec_1028 <= _zz_regVec_0;
          end
          if(_zz_1[1029]) begin
            regVec_1029 <= _zz_regVec_0;
          end
          if(_zz_1[1030]) begin
            regVec_1030 <= _zz_regVec_0;
          end
          if(_zz_1[1031]) begin
            regVec_1031 <= _zz_regVec_0;
          end
          if(_zz_1[1032]) begin
            regVec_1032 <= _zz_regVec_0;
          end
          if(_zz_1[1033]) begin
            regVec_1033 <= _zz_regVec_0;
          end
          if(_zz_1[1034]) begin
            regVec_1034 <= _zz_regVec_0;
          end
          if(_zz_1[1035]) begin
            regVec_1035 <= _zz_regVec_0;
          end
          if(_zz_1[1036]) begin
            regVec_1036 <= _zz_regVec_0;
          end
          if(_zz_1[1037]) begin
            regVec_1037 <= _zz_regVec_0;
          end
          if(_zz_1[1038]) begin
            regVec_1038 <= _zz_regVec_0;
          end
          if(_zz_1[1039]) begin
            regVec_1039 <= _zz_regVec_0;
          end
          if(_zz_1[1040]) begin
            regVec_1040 <= _zz_regVec_0;
          end
          if(_zz_1[1041]) begin
            regVec_1041 <= _zz_regVec_0;
          end
          if(_zz_1[1042]) begin
            regVec_1042 <= _zz_regVec_0;
          end
          if(_zz_1[1043]) begin
            regVec_1043 <= _zz_regVec_0;
          end
          if(_zz_1[1044]) begin
            regVec_1044 <= _zz_regVec_0;
          end
          if(_zz_1[1045]) begin
            regVec_1045 <= _zz_regVec_0;
          end
          if(_zz_1[1046]) begin
            regVec_1046 <= _zz_regVec_0;
          end
          if(_zz_1[1047]) begin
            regVec_1047 <= _zz_regVec_0;
          end
          if(_zz_1[1048]) begin
            regVec_1048 <= _zz_regVec_0;
          end
          if(_zz_1[1049]) begin
            regVec_1049 <= _zz_regVec_0;
          end
          if(_zz_1[1050]) begin
            regVec_1050 <= _zz_regVec_0;
          end
          if(_zz_1[1051]) begin
            regVec_1051 <= _zz_regVec_0;
          end
          if(_zz_1[1052]) begin
            regVec_1052 <= _zz_regVec_0;
          end
          if(_zz_1[1053]) begin
            regVec_1053 <= _zz_regVec_0;
          end
          if(_zz_1[1054]) begin
            regVec_1054 <= _zz_regVec_0;
          end
          if(_zz_1[1055]) begin
            regVec_1055 <= _zz_regVec_0;
          end
          if(_zz_1[1056]) begin
            regVec_1056 <= _zz_regVec_0;
          end
          if(_zz_1[1057]) begin
            regVec_1057 <= _zz_regVec_0;
          end
          if(_zz_1[1058]) begin
            regVec_1058 <= _zz_regVec_0;
          end
          if(_zz_1[1059]) begin
            regVec_1059 <= _zz_regVec_0;
          end
          if(_zz_1[1060]) begin
            regVec_1060 <= _zz_regVec_0;
          end
          if(_zz_1[1061]) begin
            regVec_1061 <= _zz_regVec_0;
          end
          if(_zz_1[1062]) begin
            regVec_1062 <= _zz_regVec_0;
          end
          if(_zz_1[1063]) begin
            regVec_1063 <= _zz_regVec_0;
          end
          if(_zz_1[1064]) begin
            regVec_1064 <= _zz_regVec_0;
          end
          if(_zz_1[1065]) begin
            regVec_1065 <= _zz_regVec_0;
          end
          if(_zz_1[1066]) begin
            regVec_1066 <= _zz_regVec_0;
          end
          if(_zz_1[1067]) begin
            regVec_1067 <= _zz_regVec_0;
          end
          if(_zz_1[1068]) begin
            regVec_1068 <= _zz_regVec_0;
          end
          if(_zz_1[1069]) begin
            regVec_1069 <= _zz_regVec_0;
          end
          if(_zz_1[1070]) begin
            regVec_1070 <= _zz_regVec_0;
          end
          if(_zz_1[1071]) begin
            regVec_1071 <= _zz_regVec_0;
          end
          if(_zz_1[1072]) begin
            regVec_1072 <= _zz_regVec_0;
          end
          if(_zz_1[1073]) begin
            regVec_1073 <= _zz_regVec_0;
          end
          if(_zz_1[1074]) begin
            regVec_1074 <= _zz_regVec_0;
          end
          if(_zz_1[1075]) begin
            regVec_1075 <= _zz_regVec_0;
          end
          if(_zz_1[1076]) begin
            regVec_1076 <= _zz_regVec_0;
          end
          if(_zz_1[1077]) begin
            regVec_1077 <= _zz_regVec_0;
          end
          if(_zz_1[1078]) begin
            regVec_1078 <= _zz_regVec_0;
          end
          if(_zz_1[1079]) begin
            regVec_1079 <= _zz_regVec_0;
          end
          if(_zz_1[1080]) begin
            regVec_1080 <= _zz_regVec_0;
          end
          if(_zz_1[1081]) begin
            regVec_1081 <= _zz_regVec_0;
          end
          if(_zz_1[1082]) begin
            regVec_1082 <= _zz_regVec_0;
          end
          if(_zz_1[1083]) begin
            regVec_1083 <= _zz_regVec_0;
          end
          if(_zz_1[1084]) begin
            regVec_1084 <= _zz_regVec_0;
          end
          if(_zz_1[1085]) begin
            regVec_1085 <= _zz_regVec_0;
          end
          if(_zz_1[1086]) begin
            regVec_1086 <= _zz_regVec_0;
          end
          if(_zz_1[1087]) begin
            regVec_1087 <= _zz_regVec_0;
          end
          if(_zz_1[1088]) begin
            regVec_1088 <= _zz_regVec_0;
          end
          if(_zz_1[1089]) begin
            regVec_1089 <= _zz_regVec_0;
          end
          if(_zz_1[1090]) begin
            regVec_1090 <= _zz_regVec_0;
          end
          if(_zz_1[1091]) begin
            regVec_1091 <= _zz_regVec_0;
          end
          if(_zz_1[1092]) begin
            regVec_1092 <= _zz_regVec_0;
          end
          if(_zz_1[1093]) begin
            regVec_1093 <= _zz_regVec_0;
          end
          if(_zz_1[1094]) begin
            regVec_1094 <= _zz_regVec_0;
          end
          if(_zz_1[1095]) begin
            regVec_1095 <= _zz_regVec_0;
          end
          if(_zz_1[1096]) begin
            regVec_1096 <= _zz_regVec_0;
          end
          if(_zz_1[1097]) begin
            regVec_1097 <= _zz_regVec_0;
          end
          if(_zz_1[1098]) begin
            regVec_1098 <= _zz_regVec_0;
          end
          if(_zz_1[1099]) begin
            regVec_1099 <= _zz_regVec_0;
          end
          if(_zz_1[1100]) begin
            regVec_1100 <= _zz_regVec_0;
          end
          if(_zz_1[1101]) begin
            regVec_1101 <= _zz_regVec_0;
          end
          if(_zz_1[1102]) begin
            regVec_1102 <= _zz_regVec_0;
          end
          if(_zz_1[1103]) begin
            regVec_1103 <= _zz_regVec_0;
          end
          if(_zz_1[1104]) begin
            regVec_1104 <= _zz_regVec_0;
          end
          if(_zz_1[1105]) begin
            regVec_1105 <= _zz_regVec_0;
          end
          if(_zz_1[1106]) begin
            regVec_1106 <= _zz_regVec_0;
          end
          if(_zz_1[1107]) begin
            regVec_1107 <= _zz_regVec_0;
          end
          if(_zz_1[1108]) begin
            regVec_1108 <= _zz_regVec_0;
          end
          if(_zz_1[1109]) begin
            regVec_1109 <= _zz_regVec_0;
          end
          if(_zz_1[1110]) begin
            regVec_1110 <= _zz_regVec_0;
          end
          if(_zz_1[1111]) begin
            regVec_1111 <= _zz_regVec_0;
          end
          if(_zz_1[1112]) begin
            regVec_1112 <= _zz_regVec_0;
          end
          if(_zz_1[1113]) begin
            regVec_1113 <= _zz_regVec_0;
          end
          if(_zz_1[1114]) begin
            regVec_1114 <= _zz_regVec_0;
          end
          if(_zz_1[1115]) begin
            regVec_1115 <= _zz_regVec_0;
          end
          if(_zz_1[1116]) begin
            regVec_1116 <= _zz_regVec_0;
          end
          if(_zz_1[1117]) begin
            regVec_1117 <= _zz_regVec_0;
          end
          if(_zz_1[1118]) begin
            regVec_1118 <= _zz_regVec_0;
          end
          if(_zz_1[1119]) begin
            regVec_1119 <= _zz_regVec_0;
          end
          if(_zz_1[1120]) begin
            regVec_1120 <= _zz_regVec_0;
          end
          if(_zz_1[1121]) begin
            regVec_1121 <= _zz_regVec_0;
          end
          if(_zz_1[1122]) begin
            regVec_1122 <= _zz_regVec_0;
          end
          if(_zz_1[1123]) begin
            regVec_1123 <= _zz_regVec_0;
          end
          if(_zz_1[1124]) begin
            regVec_1124 <= _zz_regVec_0;
          end
          if(_zz_1[1125]) begin
            regVec_1125 <= _zz_regVec_0;
          end
          if(_zz_1[1126]) begin
            regVec_1126 <= _zz_regVec_0;
          end
          if(_zz_1[1127]) begin
            regVec_1127 <= _zz_regVec_0;
          end
          if(_zz_1[1128]) begin
            regVec_1128 <= _zz_regVec_0;
          end
          if(_zz_1[1129]) begin
            regVec_1129 <= _zz_regVec_0;
          end
          if(_zz_1[1130]) begin
            regVec_1130 <= _zz_regVec_0;
          end
          if(_zz_1[1131]) begin
            regVec_1131 <= _zz_regVec_0;
          end
          if(_zz_1[1132]) begin
            regVec_1132 <= _zz_regVec_0;
          end
          if(_zz_1[1133]) begin
            regVec_1133 <= _zz_regVec_0;
          end
          if(_zz_1[1134]) begin
            regVec_1134 <= _zz_regVec_0;
          end
          if(_zz_1[1135]) begin
            regVec_1135 <= _zz_regVec_0;
          end
          if(_zz_1[1136]) begin
            regVec_1136 <= _zz_regVec_0;
          end
          if(_zz_1[1137]) begin
            regVec_1137 <= _zz_regVec_0;
          end
          if(_zz_1[1138]) begin
            regVec_1138 <= _zz_regVec_0;
          end
          if(_zz_1[1139]) begin
            regVec_1139 <= _zz_regVec_0;
          end
          if(_zz_1[1140]) begin
            regVec_1140 <= _zz_regVec_0;
          end
          if(_zz_1[1141]) begin
            regVec_1141 <= _zz_regVec_0;
          end
          if(_zz_1[1142]) begin
            regVec_1142 <= _zz_regVec_0;
          end
          if(_zz_1[1143]) begin
            regVec_1143 <= _zz_regVec_0;
          end
          if(_zz_1[1144]) begin
            regVec_1144 <= _zz_regVec_0;
          end
          if(_zz_1[1145]) begin
            regVec_1145 <= _zz_regVec_0;
          end
          if(_zz_1[1146]) begin
            regVec_1146 <= _zz_regVec_0;
          end
          if(_zz_1[1147]) begin
            regVec_1147 <= _zz_regVec_0;
          end
          if(_zz_1[1148]) begin
            regVec_1148 <= _zz_regVec_0;
          end
          if(_zz_1[1149]) begin
            regVec_1149 <= _zz_regVec_0;
          end
          if(_zz_1[1150]) begin
            regVec_1150 <= _zz_regVec_0;
          end
          if(_zz_1[1151]) begin
            regVec_1151 <= _zz_regVec_0;
          end
          if(_zz_1[1152]) begin
            regVec_1152 <= _zz_regVec_0;
          end
          if(_zz_1[1153]) begin
            regVec_1153 <= _zz_regVec_0;
          end
          if(_zz_1[1154]) begin
            regVec_1154 <= _zz_regVec_0;
          end
          if(_zz_1[1155]) begin
            regVec_1155 <= _zz_regVec_0;
          end
          if(_zz_1[1156]) begin
            regVec_1156 <= _zz_regVec_0;
          end
          if(_zz_1[1157]) begin
            regVec_1157 <= _zz_regVec_0;
          end
          if(_zz_1[1158]) begin
            regVec_1158 <= _zz_regVec_0;
          end
          if(_zz_1[1159]) begin
            regVec_1159 <= _zz_regVec_0;
          end
          if(_zz_1[1160]) begin
            regVec_1160 <= _zz_regVec_0;
          end
          if(_zz_1[1161]) begin
            regVec_1161 <= _zz_regVec_0;
          end
          if(_zz_1[1162]) begin
            regVec_1162 <= _zz_regVec_0;
          end
          if(_zz_1[1163]) begin
            regVec_1163 <= _zz_regVec_0;
          end
          if(_zz_1[1164]) begin
            regVec_1164 <= _zz_regVec_0;
          end
          if(_zz_1[1165]) begin
            regVec_1165 <= _zz_regVec_0;
          end
          if(_zz_1[1166]) begin
            regVec_1166 <= _zz_regVec_0;
          end
          if(_zz_1[1167]) begin
            regVec_1167 <= _zz_regVec_0;
          end
          if(_zz_1[1168]) begin
            regVec_1168 <= _zz_regVec_0;
          end
          if(_zz_1[1169]) begin
            regVec_1169 <= _zz_regVec_0;
          end
          if(_zz_1[1170]) begin
            regVec_1170 <= _zz_regVec_0;
          end
          if(_zz_1[1171]) begin
            regVec_1171 <= _zz_regVec_0;
          end
          if(_zz_1[1172]) begin
            regVec_1172 <= _zz_regVec_0;
          end
          if(_zz_1[1173]) begin
            regVec_1173 <= _zz_regVec_0;
          end
          if(_zz_1[1174]) begin
            regVec_1174 <= _zz_regVec_0;
          end
          if(_zz_1[1175]) begin
            regVec_1175 <= _zz_regVec_0;
          end
          if(_zz_1[1176]) begin
            regVec_1176 <= _zz_regVec_0;
          end
          if(_zz_1[1177]) begin
            regVec_1177 <= _zz_regVec_0;
          end
          if(_zz_1[1178]) begin
            regVec_1178 <= _zz_regVec_0;
          end
          if(_zz_1[1179]) begin
            regVec_1179 <= _zz_regVec_0;
          end
          if(_zz_1[1180]) begin
            regVec_1180 <= _zz_regVec_0;
          end
          if(_zz_1[1181]) begin
            regVec_1181 <= _zz_regVec_0;
          end
          if(_zz_1[1182]) begin
            regVec_1182 <= _zz_regVec_0;
          end
          if(_zz_1[1183]) begin
            regVec_1183 <= _zz_regVec_0;
          end
          if(_zz_1[1184]) begin
            regVec_1184 <= _zz_regVec_0;
          end
          if(_zz_1[1185]) begin
            regVec_1185 <= _zz_regVec_0;
          end
          if(_zz_1[1186]) begin
            regVec_1186 <= _zz_regVec_0;
          end
          if(_zz_1[1187]) begin
            regVec_1187 <= _zz_regVec_0;
          end
          if(_zz_1[1188]) begin
            regVec_1188 <= _zz_regVec_0;
          end
          if(_zz_1[1189]) begin
            regVec_1189 <= _zz_regVec_0;
          end
          if(_zz_1[1190]) begin
            regVec_1190 <= _zz_regVec_0;
          end
          if(_zz_1[1191]) begin
            regVec_1191 <= _zz_regVec_0;
          end
          if(_zz_1[1192]) begin
            regVec_1192 <= _zz_regVec_0;
          end
          if(_zz_1[1193]) begin
            regVec_1193 <= _zz_regVec_0;
          end
          if(_zz_1[1194]) begin
            regVec_1194 <= _zz_regVec_0;
          end
          if(_zz_1[1195]) begin
            regVec_1195 <= _zz_regVec_0;
          end
          if(_zz_1[1196]) begin
            regVec_1196 <= _zz_regVec_0;
          end
          if(_zz_1[1197]) begin
            regVec_1197 <= _zz_regVec_0;
          end
          if(_zz_1[1198]) begin
            regVec_1198 <= _zz_regVec_0;
          end
          if(_zz_1[1199]) begin
            regVec_1199 <= _zz_regVec_0;
          end
          if(_zz_1[1200]) begin
            regVec_1200 <= _zz_regVec_0;
          end
          if(_zz_1[1201]) begin
            regVec_1201 <= _zz_regVec_0;
          end
          if(_zz_1[1202]) begin
            regVec_1202 <= _zz_regVec_0;
          end
          if(_zz_1[1203]) begin
            regVec_1203 <= _zz_regVec_0;
          end
          if(_zz_1[1204]) begin
            regVec_1204 <= _zz_regVec_0;
          end
          if(_zz_1[1205]) begin
            regVec_1205 <= _zz_regVec_0;
          end
          if(_zz_1[1206]) begin
            regVec_1206 <= _zz_regVec_0;
          end
          if(_zz_1[1207]) begin
            regVec_1207 <= _zz_regVec_0;
          end
          if(_zz_1[1208]) begin
            regVec_1208 <= _zz_regVec_0;
          end
          if(_zz_1[1209]) begin
            regVec_1209 <= _zz_regVec_0;
          end
          if(_zz_1[1210]) begin
            regVec_1210 <= _zz_regVec_0;
          end
          if(_zz_1[1211]) begin
            regVec_1211 <= _zz_regVec_0;
          end
          if(_zz_1[1212]) begin
            regVec_1212 <= _zz_regVec_0;
          end
          if(_zz_1[1213]) begin
            regVec_1213 <= _zz_regVec_0;
          end
          if(_zz_1[1214]) begin
            regVec_1214 <= _zz_regVec_0;
          end
          if(_zz_1[1215]) begin
            regVec_1215 <= _zz_regVec_0;
          end
          if(_zz_1[1216]) begin
            regVec_1216 <= _zz_regVec_0;
          end
          if(_zz_1[1217]) begin
            regVec_1217 <= _zz_regVec_0;
          end
          if(_zz_1[1218]) begin
            regVec_1218 <= _zz_regVec_0;
          end
          if(_zz_1[1219]) begin
            regVec_1219 <= _zz_regVec_0;
          end
          if(_zz_1[1220]) begin
            regVec_1220 <= _zz_regVec_0;
          end
          if(_zz_1[1221]) begin
            regVec_1221 <= _zz_regVec_0;
          end
          if(_zz_1[1222]) begin
            regVec_1222 <= _zz_regVec_0;
          end
          if(_zz_1[1223]) begin
            regVec_1223 <= _zz_regVec_0;
          end
          if(_zz_1[1224]) begin
            regVec_1224 <= _zz_regVec_0;
          end
          if(_zz_1[1225]) begin
            regVec_1225 <= _zz_regVec_0;
          end
          if(_zz_1[1226]) begin
            regVec_1226 <= _zz_regVec_0;
          end
          if(_zz_1[1227]) begin
            regVec_1227 <= _zz_regVec_0;
          end
          if(_zz_1[1228]) begin
            regVec_1228 <= _zz_regVec_0;
          end
          if(_zz_1[1229]) begin
            regVec_1229 <= _zz_regVec_0;
          end
          if(_zz_1[1230]) begin
            regVec_1230 <= _zz_regVec_0;
          end
          if(_zz_1[1231]) begin
            regVec_1231 <= _zz_regVec_0;
          end
          if(_zz_1[1232]) begin
            regVec_1232 <= _zz_regVec_0;
          end
          if(_zz_1[1233]) begin
            regVec_1233 <= _zz_regVec_0;
          end
          if(_zz_1[1234]) begin
            regVec_1234 <= _zz_regVec_0;
          end
          if(_zz_1[1235]) begin
            regVec_1235 <= _zz_regVec_0;
          end
          if(_zz_1[1236]) begin
            regVec_1236 <= _zz_regVec_0;
          end
          if(_zz_1[1237]) begin
            regVec_1237 <= _zz_regVec_0;
          end
          if(_zz_1[1238]) begin
            regVec_1238 <= _zz_regVec_0;
          end
          if(_zz_1[1239]) begin
            regVec_1239 <= _zz_regVec_0;
          end
          if(_zz_1[1240]) begin
            regVec_1240 <= _zz_regVec_0;
          end
          if(_zz_1[1241]) begin
            regVec_1241 <= _zz_regVec_0;
          end
          if(_zz_1[1242]) begin
            regVec_1242 <= _zz_regVec_0;
          end
          if(_zz_1[1243]) begin
            regVec_1243 <= _zz_regVec_0;
          end
          if(_zz_1[1244]) begin
            regVec_1244 <= _zz_regVec_0;
          end
          if(_zz_1[1245]) begin
            regVec_1245 <= _zz_regVec_0;
          end
          if(_zz_1[1246]) begin
            regVec_1246 <= _zz_regVec_0;
          end
          if(_zz_1[1247]) begin
            regVec_1247 <= _zz_regVec_0;
          end
          if(_zz_1[1248]) begin
            regVec_1248 <= _zz_regVec_0;
          end
          if(_zz_1[1249]) begin
            regVec_1249 <= _zz_regVec_0;
          end
          if(_zz_1[1250]) begin
            regVec_1250 <= _zz_regVec_0;
          end
          if(_zz_1[1251]) begin
            regVec_1251 <= _zz_regVec_0;
          end
          if(_zz_1[1252]) begin
            regVec_1252 <= _zz_regVec_0;
          end
          if(_zz_1[1253]) begin
            regVec_1253 <= _zz_regVec_0;
          end
          if(_zz_1[1254]) begin
            regVec_1254 <= _zz_regVec_0;
          end
          if(_zz_1[1255]) begin
            regVec_1255 <= _zz_regVec_0;
          end
          if(_zz_1[1256]) begin
            regVec_1256 <= _zz_regVec_0;
          end
          if(_zz_1[1257]) begin
            regVec_1257 <= _zz_regVec_0;
          end
          if(_zz_1[1258]) begin
            regVec_1258 <= _zz_regVec_0;
          end
          if(_zz_1[1259]) begin
            regVec_1259 <= _zz_regVec_0;
          end
          if(_zz_1[1260]) begin
            regVec_1260 <= _zz_regVec_0;
          end
          if(_zz_1[1261]) begin
            regVec_1261 <= _zz_regVec_0;
          end
          if(_zz_1[1262]) begin
            regVec_1262 <= _zz_regVec_0;
          end
          if(_zz_1[1263]) begin
            regVec_1263 <= _zz_regVec_0;
          end
          if(_zz_1[1264]) begin
            regVec_1264 <= _zz_regVec_0;
          end
          if(_zz_1[1265]) begin
            regVec_1265 <= _zz_regVec_0;
          end
          if(_zz_1[1266]) begin
            regVec_1266 <= _zz_regVec_0;
          end
          if(_zz_1[1267]) begin
            regVec_1267 <= _zz_regVec_0;
          end
          if(_zz_1[1268]) begin
            regVec_1268 <= _zz_regVec_0;
          end
          if(_zz_1[1269]) begin
            regVec_1269 <= _zz_regVec_0;
          end
          if(_zz_1[1270]) begin
            regVec_1270 <= _zz_regVec_0;
          end
          if(_zz_1[1271]) begin
            regVec_1271 <= _zz_regVec_0;
          end
          if(_zz_1[1272]) begin
            regVec_1272 <= _zz_regVec_0;
          end
          if(_zz_1[1273]) begin
            regVec_1273 <= _zz_regVec_0;
          end
          if(_zz_1[1274]) begin
            regVec_1274 <= _zz_regVec_0;
          end
          if(_zz_1[1275]) begin
            regVec_1275 <= _zz_regVec_0;
          end
          if(_zz_1[1276]) begin
            regVec_1276 <= _zz_regVec_0;
          end
          if(_zz_1[1277]) begin
            regVec_1277 <= _zz_regVec_0;
          end
          if(_zz_1[1278]) begin
            regVec_1278 <= _zz_regVec_0;
          end
          if(_zz_1[1279]) begin
            regVec_1279 <= _zz_regVec_0;
          end
          if(_zz_1[1280]) begin
            regVec_1280 <= _zz_regVec_0;
          end
          if(_zz_1[1281]) begin
            regVec_1281 <= _zz_regVec_0;
          end
          if(_zz_1[1282]) begin
            regVec_1282 <= _zz_regVec_0;
          end
          if(_zz_1[1283]) begin
            regVec_1283 <= _zz_regVec_0;
          end
          if(_zz_1[1284]) begin
            regVec_1284 <= _zz_regVec_0;
          end
          if(_zz_1[1285]) begin
            regVec_1285 <= _zz_regVec_0;
          end
          if(_zz_1[1286]) begin
            regVec_1286 <= _zz_regVec_0;
          end
          if(_zz_1[1287]) begin
            regVec_1287 <= _zz_regVec_0;
          end
          if(_zz_1[1288]) begin
            regVec_1288 <= _zz_regVec_0;
          end
          if(_zz_1[1289]) begin
            regVec_1289 <= _zz_regVec_0;
          end
          if(_zz_1[1290]) begin
            regVec_1290 <= _zz_regVec_0;
          end
          if(_zz_1[1291]) begin
            regVec_1291 <= _zz_regVec_0;
          end
          if(_zz_1[1292]) begin
            regVec_1292 <= _zz_regVec_0;
          end
          if(_zz_1[1293]) begin
            regVec_1293 <= _zz_regVec_0;
          end
          if(_zz_1[1294]) begin
            regVec_1294 <= _zz_regVec_0;
          end
          if(_zz_1[1295]) begin
            regVec_1295 <= _zz_regVec_0;
          end
          if(_zz_1[1296]) begin
            regVec_1296 <= _zz_regVec_0;
          end
          if(_zz_1[1297]) begin
            regVec_1297 <= _zz_regVec_0;
          end
          if(_zz_1[1298]) begin
            regVec_1298 <= _zz_regVec_0;
          end
          if(_zz_1[1299]) begin
            regVec_1299 <= _zz_regVec_0;
          end
          if(_zz_1[1300]) begin
            regVec_1300 <= _zz_regVec_0;
          end
          if(_zz_1[1301]) begin
            regVec_1301 <= _zz_regVec_0;
          end
          if(_zz_1[1302]) begin
            regVec_1302 <= _zz_regVec_0;
          end
          if(_zz_1[1303]) begin
            regVec_1303 <= _zz_regVec_0;
          end
          if(_zz_1[1304]) begin
            regVec_1304 <= _zz_regVec_0;
          end
          if(_zz_1[1305]) begin
            regVec_1305 <= _zz_regVec_0;
          end
          if(_zz_1[1306]) begin
            regVec_1306 <= _zz_regVec_0;
          end
          if(_zz_1[1307]) begin
            regVec_1307 <= _zz_regVec_0;
          end
          if(_zz_1[1308]) begin
            regVec_1308 <= _zz_regVec_0;
          end
          if(_zz_1[1309]) begin
            regVec_1309 <= _zz_regVec_0;
          end
          if(_zz_1[1310]) begin
            regVec_1310 <= _zz_regVec_0;
          end
          if(_zz_1[1311]) begin
            regVec_1311 <= _zz_regVec_0;
          end
          if(_zz_1[1312]) begin
            regVec_1312 <= _zz_regVec_0;
          end
          if(_zz_1[1313]) begin
            regVec_1313 <= _zz_regVec_0;
          end
          if(_zz_1[1314]) begin
            regVec_1314 <= _zz_regVec_0;
          end
          if(_zz_1[1315]) begin
            regVec_1315 <= _zz_regVec_0;
          end
          if(_zz_1[1316]) begin
            regVec_1316 <= _zz_regVec_0;
          end
          if(_zz_1[1317]) begin
            regVec_1317 <= _zz_regVec_0;
          end
          if(_zz_1[1318]) begin
            regVec_1318 <= _zz_regVec_0;
          end
          if(_zz_1[1319]) begin
            regVec_1319 <= _zz_regVec_0;
          end
          if(_zz_1[1320]) begin
            regVec_1320 <= _zz_regVec_0;
          end
          if(_zz_1[1321]) begin
            regVec_1321 <= _zz_regVec_0;
          end
          if(_zz_1[1322]) begin
            regVec_1322 <= _zz_regVec_0;
          end
          if(_zz_1[1323]) begin
            regVec_1323 <= _zz_regVec_0;
          end
          if(_zz_1[1324]) begin
            regVec_1324 <= _zz_regVec_0;
          end
          if(_zz_1[1325]) begin
            regVec_1325 <= _zz_regVec_0;
          end
          if(_zz_1[1326]) begin
            regVec_1326 <= _zz_regVec_0;
          end
          if(_zz_1[1327]) begin
            regVec_1327 <= _zz_regVec_0;
          end
          if(_zz_1[1328]) begin
            regVec_1328 <= _zz_regVec_0;
          end
          if(_zz_1[1329]) begin
            regVec_1329 <= _zz_regVec_0;
          end
          if(_zz_1[1330]) begin
            regVec_1330 <= _zz_regVec_0;
          end
          if(_zz_1[1331]) begin
            regVec_1331 <= _zz_regVec_0;
          end
          if(_zz_1[1332]) begin
            regVec_1332 <= _zz_regVec_0;
          end
          if(_zz_1[1333]) begin
            regVec_1333 <= _zz_regVec_0;
          end
          if(_zz_1[1334]) begin
            regVec_1334 <= _zz_regVec_0;
          end
          if(_zz_1[1335]) begin
            regVec_1335 <= _zz_regVec_0;
          end
          if(_zz_1[1336]) begin
            regVec_1336 <= _zz_regVec_0;
          end
          if(_zz_1[1337]) begin
            regVec_1337 <= _zz_regVec_0;
          end
          if(_zz_1[1338]) begin
            regVec_1338 <= _zz_regVec_0;
          end
          if(_zz_1[1339]) begin
            regVec_1339 <= _zz_regVec_0;
          end
          if(_zz_1[1340]) begin
            regVec_1340 <= _zz_regVec_0;
          end
          if(_zz_1[1341]) begin
            regVec_1341 <= _zz_regVec_0;
          end
          if(_zz_1[1342]) begin
            regVec_1342 <= _zz_regVec_0;
          end
          if(_zz_1[1343]) begin
            regVec_1343 <= _zz_regVec_0;
          end
          if(_zz_1[1344]) begin
            regVec_1344 <= _zz_regVec_0;
          end
          if(_zz_1[1345]) begin
            regVec_1345 <= _zz_regVec_0;
          end
          if(_zz_1[1346]) begin
            regVec_1346 <= _zz_regVec_0;
          end
          if(_zz_1[1347]) begin
            regVec_1347 <= _zz_regVec_0;
          end
          if(_zz_1[1348]) begin
            regVec_1348 <= _zz_regVec_0;
          end
          if(_zz_1[1349]) begin
            regVec_1349 <= _zz_regVec_0;
          end
          if(_zz_1[1350]) begin
            regVec_1350 <= _zz_regVec_0;
          end
          if(_zz_1[1351]) begin
            regVec_1351 <= _zz_regVec_0;
          end
          if(_zz_1[1352]) begin
            regVec_1352 <= _zz_regVec_0;
          end
          if(_zz_1[1353]) begin
            regVec_1353 <= _zz_regVec_0;
          end
          if(_zz_1[1354]) begin
            regVec_1354 <= _zz_regVec_0;
          end
          if(_zz_1[1355]) begin
            regVec_1355 <= _zz_regVec_0;
          end
          if(_zz_1[1356]) begin
            regVec_1356 <= _zz_regVec_0;
          end
          if(_zz_1[1357]) begin
            regVec_1357 <= _zz_regVec_0;
          end
          if(_zz_1[1358]) begin
            regVec_1358 <= _zz_regVec_0;
          end
          if(_zz_1[1359]) begin
            regVec_1359 <= _zz_regVec_0;
          end
          if(_zz_1[1360]) begin
            regVec_1360 <= _zz_regVec_0;
          end
          if(_zz_1[1361]) begin
            regVec_1361 <= _zz_regVec_0;
          end
          if(_zz_1[1362]) begin
            regVec_1362 <= _zz_regVec_0;
          end
          if(_zz_1[1363]) begin
            regVec_1363 <= _zz_regVec_0;
          end
          if(_zz_1[1364]) begin
            regVec_1364 <= _zz_regVec_0;
          end
          if(_zz_1[1365]) begin
            regVec_1365 <= _zz_regVec_0;
          end
          if(_zz_1[1366]) begin
            regVec_1366 <= _zz_regVec_0;
          end
          if(_zz_1[1367]) begin
            regVec_1367 <= _zz_regVec_0;
          end
          if(_zz_1[1368]) begin
            regVec_1368 <= _zz_regVec_0;
          end
          if(_zz_1[1369]) begin
            regVec_1369 <= _zz_regVec_0;
          end
          if(_zz_1[1370]) begin
            regVec_1370 <= _zz_regVec_0;
          end
          if(_zz_1[1371]) begin
            regVec_1371 <= _zz_regVec_0;
          end
          if(_zz_1[1372]) begin
            regVec_1372 <= _zz_regVec_0;
          end
          if(_zz_1[1373]) begin
            regVec_1373 <= _zz_regVec_0;
          end
          if(_zz_1[1374]) begin
            regVec_1374 <= _zz_regVec_0;
          end
          if(_zz_1[1375]) begin
            regVec_1375 <= _zz_regVec_0;
          end
          if(_zz_1[1376]) begin
            regVec_1376 <= _zz_regVec_0;
          end
          if(_zz_1[1377]) begin
            regVec_1377 <= _zz_regVec_0;
          end
          if(_zz_1[1378]) begin
            regVec_1378 <= _zz_regVec_0;
          end
          if(_zz_1[1379]) begin
            regVec_1379 <= _zz_regVec_0;
          end
          if(_zz_1[1380]) begin
            regVec_1380 <= _zz_regVec_0;
          end
          if(_zz_1[1381]) begin
            regVec_1381 <= _zz_regVec_0;
          end
          if(_zz_1[1382]) begin
            regVec_1382 <= _zz_regVec_0;
          end
          if(_zz_1[1383]) begin
            regVec_1383 <= _zz_regVec_0;
          end
          if(_zz_1[1384]) begin
            regVec_1384 <= _zz_regVec_0;
          end
          if(_zz_1[1385]) begin
            regVec_1385 <= _zz_regVec_0;
          end
          if(_zz_1[1386]) begin
            regVec_1386 <= _zz_regVec_0;
          end
          if(_zz_1[1387]) begin
            regVec_1387 <= _zz_regVec_0;
          end
          if(_zz_1[1388]) begin
            regVec_1388 <= _zz_regVec_0;
          end
          if(_zz_1[1389]) begin
            regVec_1389 <= _zz_regVec_0;
          end
          if(_zz_1[1390]) begin
            regVec_1390 <= _zz_regVec_0;
          end
          if(_zz_1[1391]) begin
            regVec_1391 <= _zz_regVec_0;
          end
          if(_zz_1[1392]) begin
            regVec_1392 <= _zz_regVec_0;
          end
          if(_zz_1[1393]) begin
            regVec_1393 <= _zz_regVec_0;
          end
          if(_zz_1[1394]) begin
            regVec_1394 <= _zz_regVec_0;
          end
          if(_zz_1[1395]) begin
            regVec_1395 <= _zz_regVec_0;
          end
          if(_zz_1[1396]) begin
            regVec_1396 <= _zz_regVec_0;
          end
          if(_zz_1[1397]) begin
            regVec_1397 <= _zz_regVec_0;
          end
          if(_zz_1[1398]) begin
            regVec_1398 <= _zz_regVec_0;
          end
          if(_zz_1[1399]) begin
            regVec_1399 <= _zz_regVec_0;
          end
          if(_zz_1[1400]) begin
            regVec_1400 <= _zz_regVec_0;
          end
          if(_zz_1[1401]) begin
            regVec_1401 <= _zz_regVec_0;
          end
          if(_zz_1[1402]) begin
            regVec_1402 <= _zz_regVec_0;
          end
          if(_zz_1[1403]) begin
            regVec_1403 <= _zz_regVec_0;
          end
          if(_zz_1[1404]) begin
            regVec_1404 <= _zz_regVec_0;
          end
          if(_zz_1[1405]) begin
            regVec_1405 <= _zz_regVec_0;
          end
          if(_zz_1[1406]) begin
            regVec_1406 <= _zz_regVec_0;
          end
          if(_zz_1[1407]) begin
            regVec_1407 <= _zz_regVec_0;
          end
          if(_zz_1[1408]) begin
            regVec_1408 <= _zz_regVec_0;
          end
          if(_zz_1[1409]) begin
            regVec_1409 <= _zz_regVec_0;
          end
          if(_zz_1[1410]) begin
            regVec_1410 <= _zz_regVec_0;
          end
          if(_zz_1[1411]) begin
            regVec_1411 <= _zz_regVec_0;
          end
          if(_zz_1[1412]) begin
            regVec_1412 <= _zz_regVec_0;
          end
          if(_zz_1[1413]) begin
            regVec_1413 <= _zz_regVec_0;
          end
          if(_zz_1[1414]) begin
            regVec_1414 <= _zz_regVec_0;
          end
          if(_zz_1[1415]) begin
            regVec_1415 <= _zz_regVec_0;
          end
          if(_zz_1[1416]) begin
            regVec_1416 <= _zz_regVec_0;
          end
          if(_zz_1[1417]) begin
            regVec_1417 <= _zz_regVec_0;
          end
          if(_zz_1[1418]) begin
            regVec_1418 <= _zz_regVec_0;
          end
          if(_zz_1[1419]) begin
            regVec_1419 <= _zz_regVec_0;
          end
          if(_zz_1[1420]) begin
            regVec_1420 <= _zz_regVec_0;
          end
          if(_zz_1[1421]) begin
            regVec_1421 <= _zz_regVec_0;
          end
          if(_zz_1[1422]) begin
            regVec_1422 <= _zz_regVec_0;
          end
          if(_zz_1[1423]) begin
            regVec_1423 <= _zz_regVec_0;
          end
          if(_zz_1[1424]) begin
            regVec_1424 <= _zz_regVec_0;
          end
          if(_zz_1[1425]) begin
            regVec_1425 <= _zz_regVec_0;
          end
          if(_zz_1[1426]) begin
            regVec_1426 <= _zz_regVec_0;
          end
          if(_zz_1[1427]) begin
            regVec_1427 <= _zz_regVec_0;
          end
          if(_zz_1[1428]) begin
            regVec_1428 <= _zz_regVec_0;
          end
          if(_zz_1[1429]) begin
            regVec_1429 <= _zz_regVec_0;
          end
          if(_zz_1[1430]) begin
            regVec_1430 <= _zz_regVec_0;
          end
          if(_zz_1[1431]) begin
            regVec_1431 <= _zz_regVec_0;
          end
          if(_zz_1[1432]) begin
            regVec_1432 <= _zz_regVec_0;
          end
          if(_zz_1[1433]) begin
            regVec_1433 <= _zz_regVec_0;
          end
          if(_zz_1[1434]) begin
            regVec_1434 <= _zz_regVec_0;
          end
          if(_zz_1[1435]) begin
            regVec_1435 <= _zz_regVec_0;
          end
          if(_zz_1[1436]) begin
            regVec_1436 <= _zz_regVec_0;
          end
          if(_zz_1[1437]) begin
            regVec_1437 <= _zz_regVec_0;
          end
          if(_zz_1[1438]) begin
            regVec_1438 <= _zz_regVec_0;
          end
          if(_zz_1[1439]) begin
            regVec_1439 <= _zz_regVec_0;
          end
          if(_zz_1[1440]) begin
            regVec_1440 <= _zz_regVec_0;
          end
          if(_zz_1[1441]) begin
            regVec_1441 <= _zz_regVec_0;
          end
          if(_zz_1[1442]) begin
            regVec_1442 <= _zz_regVec_0;
          end
          if(_zz_1[1443]) begin
            regVec_1443 <= _zz_regVec_0;
          end
          if(_zz_1[1444]) begin
            regVec_1444 <= _zz_regVec_0;
          end
          if(_zz_1[1445]) begin
            regVec_1445 <= _zz_regVec_0;
          end
          if(_zz_1[1446]) begin
            regVec_1446 <= _zz_regVec_0;
          end
          if(_zz_1[1447]) begin
            regVec_1447 <= _zz_regVec_0;
          end
          if(_zz_1[1448]) begin
            regVec_1448 <= _zz_regVec_0;
          end
          if(_zz_1[1449]) begin
            regVec_1449 <= _zz_regVec_0;
          end
          if(_zz_1[1450]) begin
            regVec_1450 <= _zz_regVec_0;
          end
          if(_zz_1[1451]) begin
            regVec_1451 <= _zz_regVec_0;
          end
          if(_zz_1[1452]) begin
            regVec_1452 <= _zz_regVec_0;
          end
          if(_zz_1[1453]) begin
            regVec_1453 <= _zz_regVec_0;
          end
          if(_zz_1[1454]) begin
            regVec_1454 <= _zz_regVec_0;
          end
          if(_zz_1[1455]) begin
            regVec_1455 <= _zz_regVec_0;
          end
          if(_zz_1[1456]) begin
            regVec_1456 <= _zz_regVec_0;
          end
          if(_zz_1[1457]) begin
            regVec_1457 <= _zz_regVec_0;
          end
          if(_zz_1[1458]) begin
            regVec_1458 <= _zz_regVec_0;
          end
          if(_zz_1[1459]) begin
            regVec_1459 <= _zz_regVec_0;
          end
          if(_zz_1[1460]) begin
            regVec_1460 <= _zz_regVec_0;
          end
          if(_zz_1[1461]) begin
            regVec_1461 <= _zz_regVec_0;
          end
          if(_zz_1[1462]) begin
            regVec_1462 <= _zz_regVec_0;
          end
          if(_zz_1[1463]) begin
            regVec_1463 <= _zz_regVec_0;
          end
          if(_zz_1[1464]) begin
            regVec_1464 <= _zz_regVec_0;
          end
          if(_zz_1[1465]) begin
            regVec_1465 <= _zz_regVec_0;
          end
          if(_zz_1[1466]) begin
            regVec_1466 <= _zz_regVec_0;
          end
          if(_zz_1[1467]) begin
            regVec_1467 <= _zz_regVec_0;
          end
          if(_zz_1[1468]) begin
            regVec_1468 <= _zz_regVec_0;
          end
          if(_zz_1[1469]) begin
            regVec_1469 <= _zz_regVec_0;
          end
          if(_zz_1[1470]) begin
            regVec_1470 <= _zz_regVec_0;
          end
          if(_zz_1[1471]) begin
            regVec_1471 <= _zz_regVec_0;
          end
          if(_zz_1[1472]) begin
            regVec_1472 <= _zz_regVec_0;
          end
          if(_zz_1[1473]) begin
            regVec_1473 <= _zz_regVec_0;
          end
          if(_zz_1[1474]) begin
            regVec_1474 <= _zz_regVec_0;
          end
          if(_zz_1[1475]) begin
            regVec_1475 <= _zz_regVec_0;
          end
          if(_zz_1[1476]) begin
            regVec_1476 <= _zz_regVec_0;
          end
          if(_zz_1[1477]) begin
            regVec_1477 <= _zz_regVec_0;
          end
          if(_zz_1[1478]) begin
            regVec_1478 <= _zz_regVec_0;
          end
          if(_zz_1[1479]) begin
            regVec_1479 <= _zz_regVec_0;
          end
          if(_zz_1[1480]) begin
            regVec_1480 <= _zz_regVec_0;
          end
          if(_zz_1[1481]) begin
            regVec_1481 <= _zz_regVec_0;
          end
          if(_zz_1[1482]) begin
            regVec_1482 <= _zz_regVec_0;
          end
          if(_zz_1[1483]) begin
            regVec_1483 <= _zz_regVec_0;
          end
          if(_zz_1[1484]) begin
            regVec_1484 <= _zz_regVec_0;
          end
          if(_zz_1[1485]) begin
            regVec_1485 <= _zz_regVec_0;
          end
          if(_zz_1[1486]) begin
            regVec_1486 <= _zz_regVec_0;
          end
          if(_zz_1[1487]) begin
            regVec_1487 <= _zz_regVec_0;
          end
          if(_zz_1[1488]) begin
            regVec_1488 <= _zz_regVec_0;
          end
          if(_zz_1[1489]) begin
            regVec_1489 <= _zz_regVec_0;
          end
          if(_zz_1[1490]) begin
            regVec_1490 <= _zz_regVec_0;
          end
          if(_zz_1[1491]) begin
            regVec_1491 <= _zz_regVec_0;
          end
          if(_zz_1[1492]) begin
            regVec_1492 <= _zz_regVec_0;
          end
          if(_zz_1[1493]) begin
            regVec_1493 <= _zz_regVec_0;
          end
          if(_zz_1[1494]) begin
            regVec_1494 <= _zz_regVec_0;
          end
          if(_zz_1[1495]) begin
            regVec_1495 <= _zz_regVec_0;
          end
          if(_zz_1[1496]) begin
            regVec_1496 <= _zz_regVec_0;
          end
          if(_zz_1[1497]) begin
            regVec_1497 <= _zz_regVec_0;
          end
          if(_zz_1[1498]) begin
            regVec_1498 <= _zz_regVec_0;
          end
          if(_zz_1[1499]) begin
            regVec_1499 <= _zz_regVec_0;
          end
          if(_zz_1[1500]) begin
            regVec_1500 <= _zz_regVec_0;
          end
          if(_zz_1[1501]) begin
            regVec_1501 <= _zz_regVec_0;
          end
          if(_zz_1[1502]) begin
            regVec_1502 <= _zz_regVec_0;
          end
          if(_zz_1[1503]) begin
            regVec_1503 <= _zz_regVec_0;
          end
          if(_zz_1[1504]) begin
            regVec_1504 <= _zz_regVec_0;
          end
          if(_zz_1[1505]) begin
            regVec_1505 <= _zz_regVec_0;
          end
          if(_zz_1[1506]) begin
            regVec_1506 <= _zz_regVec_0;
          end
          if(_zz_1[1507]) begin
            regVec_1507 <= _zz_regVec_0;
          end
          if(_zz_1[1508]) begin
            regVec_1508 <= _zz_regVec_0;
          end
          if(_zz_1[1509]) begin
            regVec_1509 <= _zz_regVec_0;
          end
          if(_zz_1[1510]) begin
            regVec_1510 <= _zz_regVec_0;
          end
          if(_zz_1[1511]) begin
            regVec_1511 <= _zz_regVec_0;
          end
          if(_zz_1[1512]) begin
            regVec_1512 <= _zz_regVec_0;
          end
          if(_zz_1[1513]) begin
            regVec_1513 <= _zz_regVec_0;
          end
          if(_zz_1[1514]) begin
            regVec_1514 <= _zz_regVec_0;
          end
          if(_zz_1[1515]) begin
            regVec_1515 <= _zz_regVec_0;
          end
          if(_zz_1[1516]) begin
            regVec_1516 <= _zz_regVec_0;
          end
          if(_zz_1[1517]) begin
            regVec_1517 <= _zz_regVec_0;
          end
          if(_zz_1[1518]) begin
            regVec_1518 <= _zz_regVec_0;
          end
          if(_zz_1[1519]) begin
            regVec_1519 <= _zz_regVec_0;
          end
          if(_zz_1[1520]) begin
            regVec_1520 <= _zz_regVec_0;
          end
          if(_zz_1[1521]) begin
            regVec_1521 <= _zz_regVec_0;
          end
          if(_zz_1[1522]) begin
            regVec_1522 <= _zz_regVec_0;
          end
          if(_zz_1[1523]) begin
            regVec_1523 <= _zz_regVec_0;
          end
          if(_zz_1[1524]) begin
            regVec_1524 <= _zz_regVec_0;
          end
          if(_zz_1[1525]) begin
            regVec_1525 <= _zz_regVec_0;
          end
          if(_zz_1[1526]) begin
            regVec_1526 <= _zz_regVec_0;
          end
          if(_zz_1[1527]) begin
            regVec_1527 <= _zz_regVec_0;
          end
          if(_zz_1[1528]) begin
            regVec_1528 <= _zz_regVec_0;
          end
          if(_zz_1[1529]) begin
            regVec_1529 <= _zz_regVec_0;
          end
          if(_zz_1[1530]) begin
            regVec_1530 <= _zz_regVec_0;
          end
          if(_zz_1[1531]) begin
            regVec_1531 <= _zz_regVec_0;
          end
          if(_zz_1[1532]) begin
            regVec_1532 <= _zz_regVec_0;
          end
          if(_zz_1[1533]) begin
            regVec_1533 <= _zz_regVec_0;
          end
          if(_zz_1[1534]) begin
            regVec_1534 <= _zz_regVec_0;
          end
          if(_zz_1[1535]) begin
            regVec_1535 <= _zz_regVec_0;
          end
          if(_zz_1[1536]) begin
            regVec_1536 <= _zz_regVec_0;
          end
          if(_zz_1[1537]) begin
            regVec_1537 <= _zz_regVec_0;
          end
          if(_zz_1[1538]) begin
            regVec_1538 <= _zz_regVec_0;
          end
          if(_zz_1[1539]) begin
            regVec_1539 <= _zz_regVec_0;
          end
          if(_zz_1[1540]) begin
            regVec_1540 <= _zz_regVec_0;
          end
          if(_zz_1[1541]) begin
            regVec_1541 <= _zz_regVec_0;
          end
          if(_zz_1[1542]) begin
            regVec_1542 <= _zz_regVec_0;
          end
          if(_zz_1[1543]) begin
            regVec_1543 <= _zz_regVec_0;
          end
          if(_zz_1[1544]) begin
            regVec_1544 <= _zz_regVec_0;
          end
          if(_zz_1[1545]) begin
            regVec_1545 <= _zz_regVec_0;
          end
          if(_zz_1[1546]) begin
            regVec_1546 <= _zz_regVec_0;
          end
          if(_zz_1[1547]) begin
            regVec_1547 <= _zz_regVec_0;
          end
          if(_zz_1[1548]) begin
            regVec_1548 <= _zz_regVec_0;
          end
          if(_zz_1[1549]) begin
            regVec_1549 <= _zz_regVec_0;
          end
          if(_zz_1[1550]) begin
            regVec_1550 <= _zz_regVec_0;
          end
          if(_zz_1[1551]) begin
            regVec_1551 <= _zz_regVec_0;
          end
          if(_zz_1[1552]) begin
            regVec_1552 <= _zz_regVec_0;
          end
          if(_zz_1[1553]) begin
            regVec_1553 <= _zz_regVec_0;
          end
          if(_zz_1[1554]) begin
            regVec_1554 <= _zz_regVec_0;
          end
          if(_zz_1[1555]) begin
            regVec_1555 <= _zz_regVec_0;
          end
          if(_zz_1[1556]) begin
            regVec_1556 <= _zz_regVec_0;
          end
          if(_zz_1[1557]) begin
            regVec_1557 <= _zz_regVec_0;
          end
          if(_zz_1[1558]) begin
            regVec_1558 <= _zz_regVec_0;
          end
          if(_zz_1[1559]) begin
            regVec_1559 <= _zz_regVec_0;
          end
          if(_zz_1[1560]) begin
            regVec_1560 <= _zz_regVec_0;
          end
          if(_zz_1[1561]) begin
            regVec_1561 <= _zz_regVec_0;
          end
          if(_zz_1[1562]) begin
            regVec_1562 <= _zz_regVec_0;
          end
          if(_zz_1[1563]) begin
            regVec_1563 <= _zz_regVec_0;
          end
          if(_zz_1[1564]) begin
            regVec_1564 <= _zz_regVec_0;
          end
          if(_zz_1[1565]) begin
            regVec_1565 <= _zz_regVec_0;
          end
          if(_zz_1[1566]) begin
            regVec_1566 <= _zz_regVec_0;
          end
          if(_zz_1[1567]) begin
            regVec_1567 <= _zz_regVec_0;
          end
          if(_zz_1[1568]) begin
            regVec_1568 <= _zz_regVec_0;
          end
          if(_zz_1[1569]) begin
            regVec_1569 <= _zz_regVec_0;
          end
          if(_zz_1[1570]) begin
            regVec_1570 <= _zz_regVec_0;
          end
          if(_zz_1[1571]) begin
            regVec_1571 <= _zz_regVec_0;
          end
          if(_zz_1[1572]) begin
            regVec_1572 <= _zz_regVec_0;
          end
          if(_zz_1[1573]) begin
            regVec_1573 <= _zz_regVec_0;
          end
          if(_zz_1[1574]) begin
            regVec_1574 <= _zz_regVec_0;
          end
          if(_zz_1[1575]) begin
            regVec_1575 <= _zz_regVec_0;
          end
          if(_zz_1[1576]) begin
            regVec_1576 <= _zz_regVec_0;
          end
          if(_zz_1[1577]) begin
            regVec_1577 <= _zz_regVec_0;
          end
          if(_zz_1[1578]) begin
            regVec_1578 <= _zz_regVec_0;
          end
          if(_zz_1[1579]) begin
            regVec_1579 <= _zz_regVec_0;
          end
          if(_zz_1[1580]) begin
            regVec_1580 <= _zz_regVec_0;
          end
          if(_zz_1[1581]) begin
            regVec_1581 <= _zz_regVec_0;
          end
          if(_zz_1[1582]) begin
            regVec_1582 <= _zz_regVec_0;
          end
          if(_zz_1[1583]) begin
            regVec_1583 <= _zz_regVec_0;
          end
          if(_zz_1[1584]) begin
            regVec_1584 <= _zz_regVec_0;
          end
          if(_zz_1[1585]) begin
            regVec_1585 <= _zz_regVec_0;
          end
          if(_zz_1[1586]) begin
            regVec_1586 <= _zz_regVec_0;
          end
          if(_zz_1[1587]) begin
            regVec_1587 <= _zz_regVec_0;
          end
          if(_zz_1[1588]) begin
            regVec_1588 <= _zz_regVec_0;
          end
          if(_zz_1[1589]) begin
            regVec_1589 <= _zz_regVec_0;
          end
          if(_zz_1[1590]) begin
            regVec_1590 <= _zz_regVec_0;
          end
          if(_zz_1[1591]) begin
            regVec_1591 <= _zz_regVec_0;
          end
          if(_zz_1[1592]) begin
            regVec_1592 <= _zz_regVec_0;
          end
          if(_zz_1[1593]) begin
            regVec_1593 <= _zz_regVec_0;
          end
          if(_zz_1[1594]) begin
            regVec_1594 <= _zz_regVec_0;
          end
          if(_zz_1[1595]) begin
            regVec_1595 <= _zz_regVec_0;
          end
          if(_zz_1[1596]) begin
            regVec_1596 <= _zz_regVec_0;
          end
          if(_zz_1[1597]) begin
            regVec_1597 <= _zz_regVec_0;
          end
          if(_zz_1[1598]) begin
            regVec_1598 <= _zz_regVec_0;
          end
          if(_zz_1[1599]) begin
            regVec_1599 <= _zz_regVec_0;
          end
          if(_zz_1[1600]) begin
            regVec_1600 <= _zz_regVec_0;
          end
          if(_zz_1[1601]) begin
            regVec_1601 <= _zz_regVec_0;
          end
          if(_zz_1[1602]) begin
            regVec_1602 <= _zz_regVec_0;
          end
          if(_zz_1[1603]) begin
            regVec_1603 <= _zz_regVec_0;
          end
          if(_zz_1[1604]) begin
            regVec_1604 <= _zz_regVec_0;
          end
          if(_zz_1[1605]) begin
            regVec_1605 <= _zz_regVec_0;
          end
          if(_zz_1[1606]) begin
            regVec_1606 <= _zz_regVec_0;
          end
          if(_zz_1[1607]) begin
            regVec_1607 <= _zz_regVec_0;
          end
          if(_zz_1[1608]) begin
            regVec_1608 <= _zz_regVec_0;
          end
          if(_zz_1[1609]) begin
            regVec_1609 <= _zz_regVec_0;
          end
          if(_zz_1[1610]) begin
            regVec_1610 <= _zz_regVec_0;
          end
          if(_zz_1[1611]) begin
            regVec_1611 <= _zz_regVec_0;
          end
          if(_zz_1[1612]) begin
            regVec_1612 <= _zz_regVec_0;
          end
          if(_zz_1[1613]) begin
            regVec_1613 <= _zz_regVec_0;
          end
          if(_zz_1[1614]) begin
            regVec_1614 <= _zz_regVec_0;
          end
          if(_zz_1[1615]) begin
            regVec_1615 <= _zz_regVec_0;
          end
          if(_zz_1[1616]) begin
            regVec_1616 <= _zz_regVec_0;
          end
          if(_zz_1[1617]) begin
            regVec_1617 <= _zz_regVec_0;
          end
          if(_zz_1[1618]) begin
            regVec_1618 <= _zz_regVec_0;
          end
          if(_zz_1[1619]) begin
            regVec_1619 <= _zz_regVec_0;
          end
          if(_zz_1[1620]) begin
            regVec_1620 <= _zz_regVec_0;
          end
          if(_zz_1[1621]) begin
            regVec_1621 <= _zz_regVec_0;
          end
          if(_zz_1[1622]) begin
            regVec_1622 <= _zz_regVec_0;
          end
          if(_zz_1[1623]) begin
            regVec_1623 <= _zz_regVec_0;
          end
          if(_zz_1[1624]) begin
            regVec_1624 <= _zz_regVec_0;
          end
          if(_zz_1[1625]) begin
            regVec_1625 <= _zz_regVec_0;
          end
          if(_zz_1[1626]) begin
            regVec_1626 <= _zz_regVec_0;
          end
          if(_zz_1[1627]) begin
            regVec_1627 <= _zz_regVec_0;
          end
          if(_zz_1[1628]) begin
            regVec_1628 <= _zz_regVec_0;
          end
          if(_zz_1[1629]) begin
            regVec_1629 <= _zz_regVec_0;
          end
          if(_zz_1[1630]) begin
            regVec_1630 <= _zz_regVec_0;
          end
          if(_zz_1[1631]) begin
            regVec_1631 <= _zz_regVec_0;
          end
          if(_zz_1[1632]) begin
            regVec_1632 <= _zz_regVec_0;
          end
          if(_zz_1[1633]) begin
            regVec_1633 <= _zz_regVec_0;
          end
          if(_zz_1[1634]) begin
            regVec_1634 <= _zz_regVec_0;
          end
          if(_zz_1[1635]) begin
            regVec_1635 <= _zz_regVec_0;
          end
          if(_zz_1[1636]) begin
            regVec_1636 <= _zz_regVec_0;
          end
          if(_zz_1[1637]) begin
            regVec_1637 <= _zz_regVec_0;
          end
          if(_zz_1[1638]) begin
            regVec_1638 <= _zz_regVec_0;
          end
          if(_zz_1[1639]) begin
            regVec_1639 <= _zz_regVec_0;
          end
          if(_zz_1[1640]) begin
            regVec_1640 <= _zz_regVec_0;
          end
          if(_zz_1[1641]) begin
            regVec_1641 <= _zz_regVec_0;
          end
          if(_zz_1[1642]) begin
            regVec_1642 <= _zz_regVec_0;
          end
          if(_zz_1[1643]) begin
            regVec_1643 <= _zz_regVec_0;
          end
          if(_zz_1[1644]) begin
            regVec_1644 <= _zz_regVec_0;
          end
          if(_zz_1[1645]) begin
            regVec_1645 <= _zz_regVec_0;
          end
          if(_zz_1[1646]) begin
            regVec_1646 <= _zz_regVec_0;
          end
          if(_zz_1[1647]) begin
            regVec_1647 <= _zz_regVec_0;
          end
          if(_zz_1[1648]) begin
            regVec_1648 <= _zz_regVec_0;
          end
          if(_zz_1[1649]) begin
            regVec_1649 <= _zz_regVec_0;
          end
          if(_zz_1[1650]) begin
            regVec_1650 <= _zz_regVec_0;
          end
          if(_zz_1[1651]) begin
            regVec_1651 <= _zz_regVec_0;
          end
          if(_zz_1[1652]) begin
            regVec_1652 <= _zz_regVec_0;
          end
          if(_zz_1[1653]) begin
            regVec_1653 <= _zz_regVec_0;
          end
          if(_zz_1[1654]) begin
            regVec_1654 <= _zz_regVec_0;
          end
          if(_zz_1[1655]) begin
            regVec_1655 <= _zz_regVec_0;
          end
          if(_zz_1[1656]) begin
            regVec_1656 <= _zz_regVec_0;
          end
          if(_zz_1[1657]) begin
            regVec_1657 <= _zz_regVec_0;
          end
          if(_zz_1[1658]) begin
            regVec_1658 <= _zz_regVec_0;
          end
          if(_zz_1[1659]) begin
            regVec_1659 <= _zz_regVec_0;
          end
          if(_zz_1[1660]) begin
            regVec_1660 <= _zz_regVec_0;
          end
          if(_zz_1[1661]) begin
            regVec_1661 <= _zz_regVec_0;
          end
          if(_zz_1[1662]) begin
            regVec_1662 <= _zz_regVec_0;
          end
          if(_zz_1[1663]) begin
            regVec_1663 <= _zz_regVec_0;
          end
          if(_zz_1[1664]) begin
            regVec_1664 <= _zz_regVec_0;
          end
          if(_zz_1[1665]) begin
            regVec_1665 <= _zz_regVec_0;
          end
          if(_zz_1[1666]) begin
            regVec_1666 <= _zz_regVec_0;
          end
          if(_zz_1[1667]) begin
            regVec_1667 <= _zz_regVec_0;
          end
          if(_zz_1[1668]) begin
            regVec_1668 <= _zz_regVec_0;
          end
          if(_zz_1[1669]) begin
            regVec_1669 <= _zz_regVec_0;
          end
          if(_zz_1[1670]) begin
            regVec_1670 <= _zz_regVec_0;
          end
          if(_zz_1[1671]) begin
            regVec_1671 <= _zz_regVec_0;
          end
          if(_zz_1[1672]) begin
            regVec_1672 <= _zz_regVec_0;
          end
          if(_zz_1[1673]) begin
            regVec_1673 <= _zz_regVec_0;
          end
          if(_zz_1[1674]) begin
            regVec_1674 <= _zz_regVec_0;
          end
          if(_zz_1[1675]) begin
            regVec_1675 <= _zz_regVec_0;
          end
          if(_zz_1[1676]) begin
            regVec_1676 <= _zz_regVec_0;
          end
          if(_zz_1[1677]) begin
            regVec_1677 <= _zz_regVec_0;
          end
          if(_zz_1[1678]) begin
            regVec_1678 <= _zz_regVec_0;
          end
          if(_zz_1[1679]) begin
            regVec_1679 <= _zz_regVec_0;
          end
          if(_zz_1[1680]) begin
            regVec_1680 <= _zz_regVec_0;
          end
          if(_zz_1[1681]) begin
            regVec_1681 <= _zz_regVec_0;
          end
          if(_zz_1[1682]) begin
            regVec_1682 <= _zz_regVec_0;
          end
          if(_zz_1[1683]) begin
            regVec_1683 <= _zz_regVec_0;
          end
          if(_zz_1[1684]) begin
            regVec_1684 <= _zz_regVec_0;
          end
          if(_zz_1[1685]) begin
            regVec_1685 <= _zz_regVec_0;
          end
          if(_zz_1[1686]) begin
            regVec_1686 <= _zz_regVec_0;
          end
          if(_zz_1[1687]) begin
            regVec_1687 <= _zz_regVec_0;
          end
          if(_zz_1[1688]) begin
            regVec_1688 <= _zz_regVec_0;
          end
          if(_zz_1[1689]) begin
            regVec_1689 <= _zz_regVec_0;
          end
          if(_zz_1[1690]) begin
            regVec_1690 <= _zz_regVec_0;
          end
          if(_zz_1[1691]) begin
            regVec_1691 <= _zz_regVec_0;
          end
          if(_zz_1[1692]) begin
            regVec_1692 <= _zz_regVec_0;
          end
          if(_zz_1[1693]) begin
            regVec_1693 <= _zz_regVec_0;
          end
          if(_zz_1[1694]) begin
            regVec_1694 <= _zz_regVec_0;
          end
          if(_zz_1[1695]) begin
            regVec_1695 <= _zz_regVec_0;
          end
          if(_zz_1[1696]) begin
            regVec_1696 <= _zz_regVec_0;
          end
          if(_zz_1[1697]) begin
            regVec_1697 <= _zz_regVec_0;
          end
          if(_zz_1[1698]) begin
            regVec_1698 <= _zz_regVec_0;
          end
          if(_zz_1[1699]) begin
            regVec_1699 <= _zz_regVec_0;
          end
          if(_zz_1[1700]) begin
            regVec_1700 <= _zz_regVec_0;
          end
          if(_zz_1[1701]) begin
            regVec_1701 <= _zz_regVec_0;
          end
          if(_zz_1[1702]) begin
            regVec_1702 <= _zz_regVec_0;
          end
          if(_zz_1[1703]) begin
            regVec_1703 <= _zz_regVec_0;
          end
          if(_zz_1[1704]) begin
            regVec_1704 <= _zz_regVec_0;
          end
          if(_zz_1[1705]) begin
            regVec_1705 <= _zz_regVec_0;
          end
          if(_zz_1[1706]) begin
            regVec_1706 <= _zz_regVec_0;
          end
          if(_zz_1[1707]) begin
            regVec_1707 <= _zz_regVec_0;
          end
          if(_zz_1[1708]) begin
            regVec_1708 <= _zz_regVec_0;
          end
          if(_zz_1[1709]) begin
            regVec_1709 <= _zz_regVec_0;
          end
          if(_zz_1[1710]) begin
            regVec_1710 <= _zz_regVec_0;
          end
          if(_zz_1[1711]) begin
            regVec_1711 <= _zz_regVec_0;
          end
          if(_zz_1[1712]) begin
            regVec_1712 <= _zz_regVec_0;
          end
          if(_zz_1[1713]) begin
            regVec_1713 <= _zz_regVec_0;
          end
          if(_zz_1[1714]) begin
            regVec_1714 <= _zz_regVec_0;
          end
          if(_zz_1[1715]) begin
            regVec_1715 <= _zz_regVec_0;
          end
          if(_zz_1[1716]) begin
            regVec_1716 <= _zz_regVec_0;
          end
          if(_zz_1[1717]) begin
            regVec_1717 <= _zz_regVec_0;
          end
          if(_zz_1[1718]) begin
            regVec_1718 <= _zz_regVec_0;
          end
          if(_zz_1[1719]) begin
            regVec_1719 <= _zz_regVec_0;
          end
          if(_zz_1[1720]) begin
            regVec_1720 <= _zz_regVec_0;
          end
          if(_zz_1[1721]) begin
            regVec_1721 <= _zz_regVec_0;
          end
          if(_zz_1[1722]) begin
            regVec_1722 <= _zz_regVec_0;
          end
          if(_zz_1[1723]) begin
            regVec_1723 <= _zz_regVec_0;
          end
          if(_zz_1[1724]) begin
            regVec_1724 <= _zz_regVec_0;
          end
          if(_zz_1[1725]) begin
            regVec_1725 <= _zz_regVec_0;
          end
          if(_zz_1[1726]) begin
            regVec_1726 <= _zz_regVec_0;
          end
          if(_zz_1[1727]) begin
            regVec_1727 <= _zz_regVec_0;
          end
          if(_zz_1[1728]) begin
            regVec_1728 <= _zz_regVec_0;
          end
          if(_zz_1[1729]) begin
            regVec_1729 <= _zz_regVec_0;
          end
          if(_zz_1[1730]) begin
            regVec_1730 <= _zz_regVec_0;
          end
          if(_zz_1[1731]) begin
            regVec_1731 <= _zz_regVec_0;
          end
          if(_zz_1[1732]) begin
            regVec_1732 <= _zz_regVec_0;
          end
          if(_zz_1[1733]) begin
            regVec_1733 <= _zz_regVec_0;
          end
          if(_zz_1[1734]) begin
            regVec_1734 <= _zz_regVec_0;
          end
          if(_zz_1[1735]) begin
            regVec_1735 <= _zz_regVec_0;
          end
          if(_zz_1[1736]) begin
            regVec_1736 <= _zz_regVec_0;
          end
          if(_zz_1[1737]) begin
            regVec_1737 <= _zz_regVec_0;
          end
          if(_zz_1[1738]) begin
            regVec_1738 <= _zz_regVec_0;
          end
          if(_zz_1[1739]) begin
            regVec_1739 <= _zz_regVec_0;
          end
          if(_zz_1[1740]) begin
            regVec_1740 <= _zz_regVec_0;
          end
          if(_zz_1[1741]) begin
            regVec_1741 <= _zz_regVec_0;
          end
          if(_zz_1[1742]) begin
            regVec_1742 <= _zz_regVec_0;
          end
          if(_zz_1[1743]) begin
            regVec_1743 <= _zz_regVec_0;
          end
          if(_zz_1[1744]) begin
            regVec_1744 <= _zz_regVec_0;
          end
          if(_zz_1[1745]) begin
            regVec_1745 <= _zz_regVec_0;
          end
          if(_zz_1[1746]) begin
            regVec_1746 <= _zz_regVec_0;
          end
          if(_zz_1[1747]) begin
            regVec_1747 <= _zz_regVec_0;
          end
          if(_zz_1[1748]) begin
            regVec_1748 <= _zz_regVec_0;
          end
          if(_zz_1[1749]) begin
            regVec_1749 <= _zz_regVec_0;
          end
          if(_zz_1[1750]) begin
            regVec_1750 <= _zz_regVec_0;
          end
          if(_zz_1[1751]) begin
            regVec_1751 <= _zz_regVec_0;
          end
          if(_zz_1[1752]) begin
            regVec_1752 <= _zz_regVec_0;
          end
          if(_zz_1[1753]) begin
            regVec_1753 <= _zz_regVec_0;
          end
          if(_zz_1[1754]) begin
            regVec_1754 <= _zz_regVec_0;
          end
          if(_zz_1[1755]) begin
            regVec_1755 <= _zz_regVec_0;
          end
          if(_zz_1[1756]) begin
            regVec_1756 <= _zz_regVec_0;
          end
          if(_zz_1[1757]) begin
            regVec_1757 <= _zz_regVec_0;
          end
          if(_zz_1[1758]) begin
            regVec_1758 <= _zz_regVec_0;
          end
          if(_zz_1[1759]) begin
            regVec_1759 <= _zz_regVec_0;
          end
          if(_zz_1[1760]) begin
            regVec_1760 <= _zz_regVec_0;
          end
          if(_zz_1[1761]) begin
            regVec_1761 <= _zz_regVec_0;
          end
          if(_zz_1[1762]) begin
            regVec_1762 <= _zz_regVec_0;
          end
          if(_zz_1[1763]) begin
            regVec_1763 <= _zz_regVec_0;
          end
          if(_zz_1[1764]) begin
            regVec_1764 <= _zz_regVec_0;
          end
          if(_zz_1[1765]) begin
            regVec_1765 <= _zz_regVec_0;
          end
          if(_zz_1[1766]) begin
            regVec_1766 <= _zz_regVec_0;
          end
          if(_zz_1[1767]) begin
            regVec_1767 <= _zz_regVec_0;
          end
          if(_zz_1[1768]) begin
            regVec_1768 <= _zz_regVec_0;
          end
          if(_zz_1[1769]) begin
            regVec_1769 <= _zz_regVec_0;
          end
          if(_zz_1[1770]) begin
            regVec_1770 <= _zz_regVec_0;
          end
          if(_zz_1[1771]) begin
            regVec_1771 <= _zz_regVec_0;
          end
          if(_zz_1[1772]) begin
            regVec_1772 <= _zz_regVec_0;
          end
          if(_zz_1[1773]) begin
            regVec_1773 <= _zz_regVec_0;
          end
          if(_zz_1[1774]) begin
            regVec_1774 <= _zz_regVec_0;
          end
          if(_zz_1[1775]) begin
            regVec_1775 <= _zz_regVec_0;
          end
          if(_zz_1[1776]) begin
            regVec_1776 <= _zz_regVec_0;
          end
          if(_zz_1[1777]) begin
            regVec_1777 <= _zz_regVec_0;
          end
          if(_zz_1[1778]) begin
            regVec_1778 <= _zz_regVec_0;
          end
          if(_zz_1[1779]) begin
            regVec_1779 <= _zz_regVec_0;
          end
          if(_zz_1[1780]) begin
            regVec_1780 <= _zz_regVec_0;
          end
          if(_zz_1[1781]) begin
            regVec_1781 <= _zz_regVec_0;
          end
          if(_zz_1[1782]) begin
            regVec_1782 <= _zz_regVec_0;
          end
          if(_zz_1[1783]) begin
            regVec_1783 <= _zz_regVec_0;
          end
          if(_zz_1[1784]) begin
            regVec_1784 <= _zz_regVec_0;
          end
          if(_zz_1[1785]) begin
            regVec_1785 <= _zz_regVec_0;
          end
          if(_zz_1[1786]) begin
            regVec_1786 <= _zz_regVec_0;
          end
          if(_zz_1[1787]) begin
            regVec_1787 <= _zz_regVec_0;
          end
          if(_zz_1[1788]) begin
            regVec_1788 <= _zz_regVec_0;
          end
          if(_zz_1[1789]) begin
            regVec_1789 <= _zz_regVec_0;
          end
          if(_zz_1[1790]) begin
            regVec_1790 <= _zz_regVec_0;
          end
          if(_zz_1[1791]) begin
            regVec_1791 <= _zz_regVec_0;
          end
          if(_zz_1[1792]) begin
            regVec_1792 <= _zz_regVec_0;
          end
          if(_zz_1[1793]) begin
            regVec_1793 <= _zz_regVec_0;
          end
          if(_zz_1[1794]) begin
            regVec_1794 <= _zz_regVec_0;
          end
          if(_zz_1[1795]) begin
            regVec_1795 <= _zz_regVec_0;
          end
          if(_zz_1[1796]) begin
            regVec_1796 <= _zz_regVec_0;
          end
          if(_zz_1[1797]) begin
            regVec_1797 <= _zz_regVec_0;
          end
          if(_zz_1[1798]) begin
            regVec_1798 <= _zz_regVec_0;
          end
          if(_zz_1[1799]) begin
            regVec_1799 <= _zz_regVec_0;
          end
          if(_zz_1[1800]) begin
            regVec_1800 <= _zz_regVec_0;
          end
          if(_zz_1[1801]) begin
            regVec_1801 <= _zz_regVec_0;
          end
          if(_zz_1[1802]) begin
            regVec_1802 <= _zz_regVec_0;
          end
          if(_zz_1[1803]) begin
            regVec_1803 <= _zz_regVec_0;
          end
          if(_zz_1[1804]) begin
            regVec_1804 <= _zz_regVec_0;
          end
          if(_zz_1[1805]) begin
            regVec_1805 <= _zz_regVec_0;
          end
          if(_zz_1[1806]) begin
            regVec_1806 <= _zz_regVec_0;
          end
          if(_zz_1[1807]) begin
            regVec_1807 <= _zz_regVec_0;
          end
          if(_zz_1[1808]) begin
            regVec_1808 <= _zz_regVec_0;
          end
          if(_zz_1[1809]) begin
            regVec_1809 <= _zz_regVec_0;
          end
          if(_zz_1[1810]) begin
            regVec_1810 <= _zz_regVec_0;
          end
          if(_zz_1[1811]) begin
            regVec_1811 <= _zz_regVec_0;
          end
          if(_zz_1[1812]) begin
            regVec_1812 <= _zz_regVec_0;
          end
          if(_zz_1[1813]) begin
            regVec_1813 <= _zz_regVec_0;
          end
          if(_zz_1[1814]) begin
            regVec_1814 <= _zz_regVec_0;
          end
          if(_zz_1[1815]) begin
            regVec_1815 <= _zz_regVec_0;
          end
          if(_zz_1[1816]) begin
            regVec_1816 <= _zz_regVec_0;
          end
          if(_zz_1[1817]) begin
            regVec_1817 <= _zz_regVec_0;
          end
          if(_zz_1[1818]) begin
            regVec_1818 <= _zz_regVec_0;
          end
          if(_zz_1[1819]) begin
            regVec_1819 <= _zz_regVec_0;
          end
          if(_zz_1[1820]) begin
            regVec_1820 <= _zz_regVec_0;
          end
          if(_zz_1[1821]) begin
            regVec_1821 <= _zz_regVec_0;
          end
          if(_zz_1[1822]) begin
            regVec_1822 <= _zz_regVec_0;
          end
          if(_zz_1[1823]) begin
            regVec_1823 <= _zz_regVec_0;
          end
          if(_zz_1[1824]) begin
            regVec_1824 <= _zz_regVec_0;
          end
          if(_zz_1[1825]) begin
            regVec_1825 <= _zz_regVec_0;
          end
          if(_zz_1[1826]) begin
            regVec_1826 <= _zz_regVec_0;
          end
          if(_zz_1[1827]) begin
            regVec_1827 <= _zz_regVec_0;
          end
          if(_zz_1[1828]) begin
            regVec_1828 <= _zz_regVec_0;
          end
          if(_zz_1[1829]) begin
            regVec_1829 <= _zz_regVec_0;
          end
          if(_zz_1[1830]) begin
            regVec_1830 <= _zz_regVec_0;
          end
          if(_zz_1[1831]) begin
            regVec_1831 <= _zz_regVec_0;
          end
          if(_zz_1[1832]) begin
            regVec_1832 <= _zz_regVec_0;
          end
          if(_zz_1[1833]) begin
            regVec_1833 <= _zz_regVec_0;
          end
          if(_zz_1[1834]) begin
            regVec_1834 <= _zz_regVec_0;
          end
          if(_zz_1[1835]) begin
            regVec_1835 <= _zz_regVec_0;
          end
          if(_zz_1[1836]) begin
            regVec_1836 <= _zz_regVec_0;
          end
          if(_zz_1[1837]) begin
            regVec_1837 <= _zz_regVec_0;
          end
          if(_zz_1[1838]) begin
            regVec_1838 <= _zz_regVec_0;
          end
          if(_zz_1[1839]) begin
            regVec_1839 <= _zz_regVec_0;
          end
          if(_zz_1[1840]) begin
            regVec_1840 <= _zz_regVec_0;
          end
          if(_zz_1[1841]) begin
            regVec_1841 <= _zz_regVec_0;
          end
          if(_zz_1[1842]) begin
            regVec_1842 <= _zz_regVec_0;
          end
          if(_zz_1[1843]) begin
            regVec_1843 <= _zz_regVec_0;
          end
          if(_zz_1[1844]) begin
            regVec_1844 <= _zz_regVec_0;
          end
          if(_zz_1[1845]) begin
            regVec_1845 <= _zz_regVec_0;
          end
          if(_zz_1[1846]) begin
            regVec_1846 <= _zz_regVec_0;
          end
          if(_zz_1[1847]) begin
            regVec_1847 <= _zz_regVec_0;
          end
          if(_zz_1[1848]) begin
            regVec_1848 <= _zz_regVec_0;
          end
          if(_zz_1[1849]) begin
            regVec_1849 <= _zz_regVec_0;
          end
          if(_zz_1[1850]) begin
            regVec_1850 <= _zz_regVec_0;
          end
          if(_zz_1[1851]) begin
            regVec_1851 <= _zz_regVec_0;
          end
          if(_zz_1[1852]) begin
            regVec_1852 <= _zz_regVec_0;
          end
          if(_zz_1[1853]) begin
            regVec_1853 <= _zz_regVec_0;
          end
          if(_zz_1[1854]) begin
            regVec_1854 <= _zz_regVec_0;
          end
          if(_zz_1[1855]) begin
            regVec_1855 <= _zz_regVec_0;
          end
          if(_zz_1[1856]) begin
            regVec_1856 <= _zz_regVec_0;
          end
          if(_zz_1[1857]) begin
            regVec_1857 <= _zz_regVec_0;
          end
          if(_zz_1[1858]) begin
            regVec_1858 <= _zz_regVec_0;
          end
          if(_zz_1[1859]) begin
            regVec_1859 <= _zz_regVec_0;
          end
          if(_zz_1[1860]) begin
            regVec_1860 <= _zz_regVec_0;
          end
          if(_zz_1[1861]) begin
            regVec_1861 <= _zz_regVec_0;
          end
          if(_zz_1[1862]) begin
            regVec_1862 <= _zz_regVec_0;
          end
          if(_zz_1[1863]) begin
            regVec_1863 <= _zz_regVec_0;
          end
          if(_zz_1[1864]) begin
            regVec_1864 <= _zz_regVec_0;
          end
          if(_zz_1[1865]) begin
            regVec_1865 <= _zz_regVec_0;
          end
          if(_zz_1[1866]) begin
            regVec_1866 <= _zz_regVec_0;
          end
          if(_zz_1[1867]) begin
            regVec_1867 <= _zz_regVec_0;
          end
          if(_zz_1[1868]) begin
            regVec_1868 <= _zz_regVec_0;
          end
          if(_zz_1[1869]) begin
            regVec_1869 <= _zz_regVec_0;
          end
          if(_zz_1[1870]) begin
            regVec_1870 <= _zz_regVec_0;
          end
          if(_zz_1[1871]) begin
            regVec_1871 <= _zz_regVec_0;
          end
          if(_zz_1[1872]) begin
            regVec_1872 <= _zz_regVec_0;
          end
          if(_zz_1[1873]) begin
            regVec_1873 <= _zz_regVec_0;
          end
          if(_zz_1[1874]) begin
            regVec_1874 <= _zz_regVec_0;
          end
          if(_zz_1[1875]) begin
            regVec_1875 <= _zz_regVec_0;
          end
          if(_zz_1[1876]) begin
            regVec_1876 <= _zz_regVec_0;
          end
          if(_zz_1[1877]) begin
            regVec_1877 <= _zz_regVec_0;
          end
          if(_zz_1[1878]) begin
            regVec_1878 <= _zz_regVec_0;
          end
          if(_zz_1[1879]) begin
            regVec_1879 <= _zz_regVec_0;
          end
          if(_zz_1[1880]) begin
            regVec_1880 <= _zz_regVec_0;
          end
          if(_zz_1[1881]) begin
            regVec_1881 <= _zz_regVec_0;
          end
          if(_zz_1[1882]) begin
            regVec_1882 <= _zz_regVec_0;
          end
          if(_zz_1[1883]) begin
            regVec_1883 <= _zz_regVec_0;
          end
          if(_zz_1[1884]) begin
            regVec_1884 <= _zz_regVec_0;
          end
          if(_zz_1[1885]) begin
            regVec_1885 <= _zz_regVec_0;
          end
          if(_zz_1[1886]) begin
            regVec_1886 <= _zz_regVec_0;
          end
          if(_zz_1[1887]) begin
            regVec_1887 <= _zz_regVec_0;
          end
          if(_zz_1[1888]) begin
            regVec_1888 <= _zz_regVec_0;
          end
          if(_zz_1[1889]) begin
            regVec_1889 <= _zz_regVec_0;
          end
          if(_zz_1[1890]) begin
            regVec_1890 <= _zz_regVec_0;
          end
          if(_zz_1[1891]) begin
            regVec_1891 <= _zz_regVec_0;
          end
          if(_zz_1[1892]) begin
            regVec_1892 <= _zz_regVec_0;
          end
          if(_zz_1[1893]) begin
            regVec_1893 <= _zz_regVec_0;
          end
          if(_zz_1[1894]) begin
            regVec_1894 <= _zz_regVec_0;
          end
          if(_zz_1[1895]) begin
            regVec_1895 <= _zz_regVec_0;
          end
          if(_zz_1[1896]) begin
            regVec_1896 <= _zz_regVec_0;
          end
          if(_zz_1[1897]) begin
            regVec_1897 <= _zz_regVec_0;
          end
          if(_zz_1[1898]) begin
            regVec_1898 <= _zz_regVec_0;
          end
          if(_zz_1[1899]) begin
            regVec_1899 <= _zz_regVec_0;
          end
          if(_zz_1[1900]) begin
            regVec_1900 <= _zz_regVec_0;
          end
          if(_zz_1[1901]) begin
            regVec_1901 <= _zz_regVec_0;
          end
          if(_zz_1[1902]) begin
            regVec_1902 <= _zz_regVec_0;
          end
          if(_zz_1[1903]) begin
            regVec_1903 <= _zz_regVec_0;
          end
          if(_zz_1[1904]) begin
            regVec_1904 <= _zz_regVec_0;
          end
          if(_zz_1[1905]) begin
            regVec_1905 <= _zz_regVec_0;
          end
          if(_zz_1[1906]) begin
            regVec_1906 <= _zz_regVec_0;
          end
          if(_zz_1[1907]) begin
            regVec_1907 <= _zz_regVec_0;
          end
          if(_zz_1[1908]) begin
            regVec_1908 <= _zz_regVec_0;
          end
          if(_zz_1[1909]) begin
            regVec_1909 <= _zz_regVec_0;
          end
          if(_zz_1[1910]) begin
            regVec_1910 <= _zz_regVec_0;
          end
          if(_zz_1[1911]) begin
            regVec_1911 <= _zz_regVec_0;
          end
          if(_zz_1[1912]) begin
            regVec_1912 <= _zz_regVec_0;
          end
          if(_zz_1[1913]) begin
            regVec_1913 <= _zz_regVec_0;
          end
          if(_zz_1[1914]) begin
            regVec_1914 <= _zz_regVec_0;
          end
          if(_zz_1[1915]) begin
            regVec_1915 <= _zz_regVec_0;
          end
          if(_zz_1[1916]) begin
            regVec_1916 <= _zz_regVec_0;
          end
          if(_zz_1[1917]) begin
            regVec_1917 <= _zz_regVec_0;
          end
          if(_zz_1[1918]) begin
            regVec_1918 <= _zz_regVec_0;
          end
          if(_zz_1[1919]) begin
            regVec_1919 <= _zz_regVec_0;
          end
          if(_zz_1[1920]) begin
            regVec_1920 <= _zz_regVec_0;
          end
          if(_zz_1[1921]) begin
            regVec_1921 <= _zz_regVec_0;
          end
          if(_zz_1[1922]) begin
            regVec_1922 <= _zz_regVec_0;
          end
          if(_zz_1[1923]) begin
            regVec_1923 <= _zz_regVec_0;
          end
          if(_zz_1[1924]) begin
            regVec_1924 <= _zz_regVec_0;
          end
          if(_zz_1[1925]) begin
            regVec_1925 <= _zz_regVec_0;
          end
          if(_zz_1[1926]) begin
            regVec_1926 <= _zz_regVec_0;
          end
          if(_zz_1[1927]) begin
            regVec_1927 <= _zz_regVec_0;
          end
          if(_zz_1[1928]) begin
            regVec_1928 <= _zz_regVec_0;
          end
          if(_zz_1[1929]) begin
            regVec_1929 <= _zz_regVec_0;
          end
          if(_zz_1[1930]) begin
            regVec_1930 <= _zz_regVec_0;
          end
          if(_zz_1[1931]) begin
            regVec_1931 <= _zz_regVec_0;
          end
          if(_zz_1[1932]) begin
            regVec_1932 <= _zz_regVec_0;
          end
          if(_zz_1[1933]) begin
            regVec_1933 <= _zz_regVec_0;
          end
          if(_zz_1[1934]) begin
            regVec_1934 <= _zz_regVec_0;
          end
          if(_zz_1[1935]) begin
            regVec_1935 <= _zz_regVec_0;
          end
          if(_zz_1[1936]) begin
            regVec_1936 <= _zz_regVec_0;
          end
          if(_zz_1[1937]) begin
            regVec_1937 <= _zz_regVec_0;
          end
          if(_zz_1[1938]) begin
            regVec_1938 <= _zz_regVec_0;
          end
          if(_zz_1[1939]) begin
            regVec_1939 <= _zz_regVec_0;
          end
          if(_zz_1[1940]) begin
            regVec_1940 <= _zz_regVec_0;
          end
          if(_zz_1[1941]) begin
            regVec_1941 <= _zz_regVec_0;
          end
          if(_zz_1[1942]) begin
            regVec_1942 <= _zz_regVec_0;
          end
          if(_zz_1[1943]) begin
            regVec_1943 <= _zz_regVec_0;
          end
          if(_zz_1[1944]) begin
            regVec_1944 <= _zz_regVec_0;
          end
          if(_zz_1[1945]) begin
            regVec_1945 <= _zz_regVec_0;
          end
          if(_zz_1[1946]) begin
            regVec_1946 <= _zz_regVec_0;
          end
          if(_zz_1[1947]) begin
            regVec_1947 <= _zz_regVec_0;
          end
          if(_zz_1[1948]) begin
            regVec_1948 <= _zz_regVec_0;
          end
          if(_zz_1[1949]) begin
            regVec_1949 <= _zz_regVec_0;
          end
          if(_zz_1[1950]) begin
            regVec_1950 <= _zz_regVec_0;
          end
          if(_zz_1[1951]) begin
            regVec_1951 <= _zz_regVec_0;
          end
          if(_zz_1[1952]) begin
            regVec_1952 <= _zz_regVec_0;
          end
          if(_zz_1[1953]) begin
            regVec_1953 <= _zz_regVec_0;
          end
          if(_zz_1[1954]) begin
            regVec_1954 <= _zz_regVec_0;
          end
          if(_zz_1[1955]) begin
            regVec_1955 <= _zz_regVec_0;
          end
          if(_zz_1[1956]) begin
            regVec_1956 <= _zz_regVec_0;
          end
          if(_zz_1[1957]) begin
            regVec_1957 <= _zz_regVec_0;
          end
          if(_zz_1[1958]) begin
            regVec_1958 <= _zz_regVec_0;
          end
          if(_zz_1[1959]) begin
            regVec_1959 <= _zz_regVec_0;
          end
          if(_zz_1[1960]) begin
            regVec_1960 <= _zz_regVec_0;
          end
          if(_zz_1[1961]) begin
            regVec_1961 <= _zz_regVec_0;
          end
          if(_zz_1[1962]) begin
            regVec_1962 <= _zz_regVec_0;
          end
          if(_zz_1[1963]) begin
            regVec_1963 <= _zz_regVec_0;
          end
          if(_zz_1[1964]) begin
            regVec_1964 <= _zz_regVec_0;
          end
          if(_zz_1[1965]) begin
            regVec_1965 <= _zz_regVec_0;
          end
          if(_zz_1[1966]) begin
            regVec_1966 <= _zz_regVec_0;
          end
          if(_zz_1[1967]) begin
            regVec_1967 <= _zz_regVec_0;
          end
          if(_zz_1[1968]) begin
            regVec_1968 <= _zz_regVec_0;
          end
          if(_zz_1[1969]) begin
            regVec_1969 <= _zz_regVec_0;
          end
          if(_zz_1[1970]) begin
            regVec_1970 <= _zz_regVec_0;
          end
          if(_zz_1[1971]) begin
            regVec_1971 <= _zz_regVec_0;
          end
          if(_zz_1[1972]) begin
            regVec_1972 <= _zz_regVec_0;
          end
          if(_zz_1[1973]) begin
            regVec_1973 <= _zz_regVec_0;
          end
          if(_zz_1[1974]) begin
            regVec_1974 <= _zz_regVec_0;
          end
          if(_zz_1[1975]) begin
            regVec_1975 <= _zz_regVec_0;
          end
          if(_zz_1[1976]) begin
            regVec_1976 <= _zz_regVec_0;
          end
          if(_zz_1[1977]) begin
            regVec_1977 <= _zz_regVec_0;
          end
          if(_zz_1[1978]) begin
            regVec_1978 <= _zz_regVec_0;
          end
          if(_zz_1[1979]) begin
            regVec_1979 <= _zz_regVec_0;
          end
          if(_zz_1[1980]) begin
            regVec_1980 <= _zz_regVec_0;
          end
          if(_zz_1[1981]) begin
            regVec_1981 <= _zz_regVec_0;
          end
          if(_zz_1[1982]) begin
            regVec_1982 <= _zz_regVec_0;
          end
          if(_zz_1[1983]) begin
            regVec_1983 <= _zz_regVec_0;
          end
          if(_zz_1[1984]) begin
            regVec_1984 <= _zz_regVec_0;
          end
          if(_zz_1[1985]) begin
            regVec_1985 <= _zz_regVec_0;
          end
          if(_zz_1[1986]) begin
            regVec_1986 <= _zz_regVec_0;
          end
          if(_zz_1[1987]) begin
            regVec_1987 <= _zz_regVec_0;
          end
          if(_zz_1[1988]) begin
            regVec_1988 <= _zz_regVec_0;
          end
          if(_zz_1[1989]) begin
            regVec_1989 <= _zz_regVec_0;
          end
          if(_zz_1[1990]) begin
            regVec_1990 <= _zz_regVec_0;
          end
          if(_zz_1[1991]) begin
            regVec_1991 <= _zz_regVec_0;
          end
          if(_zz_1[1992]) begin
            regVec_1992 <= _zz_regVec_0;
          end
          if(_zz_1[1993]) begin
            regVec_1993 <= _zz_regVec_0;
          end
          if(_zz_1[1994]) begin
            regVec_1994 <= _zz_regVec_0;
          end
          if(_zz_1[1995]) begin
            regVec_1995 <= _zz_regVec_0;
          end
          if(_zz_1[1996]) begin
            regVec_1996 <= _zz_regVec_0;
          end
          if(_zz_1[1997]) begin
            regVec_1997 <= _zz_regVec_0;
          end
          if(_zz_1[1998]) begin
            regVec_1998 <= _zz_regVec_0;
          end
          if(_zz_1[1999]) begin
            regVec_1999 <= _zz_regVec_0;
          end
          if(_zz_1[2000]) begin
            regVec_2000 <= _zz_regVec_0;
          end
          if(_zz_1[2001]) begin
            regVec_2001 <= _zz_regVec_0;
          end
          if(_zz_1[2002]) begin
            regVec_2002 <= _zz_regVec_0;
          end
          if(_zz_1[2003]) begin
            regVec_2003 <= _zz_regVec_0;
          end
          if(_zz_1[2004]) begin
            regVec_2004 <= _zz_regVec_0;
          end
          if(_zz_1[2005]) begin
            regVec_2005 <= _zz_regVec_0;
          end
          if(_zz_1[2006]) begin
            regVec_2006 <= _zz_regVec_0;
          end
          if(_zz_1[2007]) begin
            regVec_2007 <= _zz_regVec_0;
          end
          if(_zz_1[2008]) begin
            regVec_2008 <= _zz_regVec_0;
          end
          if(_zz_1[2009]) begin
            regVec_2009 <= _zz_regVec_0;
          end
          if(_zz_1[2010]) begin
            regVec_2010 <= _zz_regVec_0;
          end
          if(_zz_1[2011]) begin
            regVec_2011 <= _zz_regVec_0;
          end
          if(_zz_1[2012]) begin
            regVec_2012 <= _zz_regVec_0;
          end
          if(_zz_1[2013]) begin
            regVec_2013 <= _zz_regVec_0;
          end
          if(_zz_1[2014]) begin
            regVec_2014 <= _zz_regVec_0;
          end
          if(_zz_1[2015]) begin
            regVec_2015 <= _zz_regVec_0;
          end
          if(_zz_1[2016]) begin
            regVec_2016 <= _zz_regVec_0;
          end
          if(_zz_1[2017]) begin
            regVec_2017 <= _zz_regVec_0;
          end
          if(_zz_1[2018]) begin
            regVec_2018 <= _zz_regVec_0;
          end
          if(_zz_1[2019]) begin
            regVec_2019 <= _zz_regVec_0;
          end
          if(_zz_1[2020]) begin
            regVec_2020 <= _zz_regVec_0;
          end
          if(_zz_1[2021]) begin
            regVec_2021 <= _zz_regVec_0;
          end
          if(_zz_1[2022]) begin
            regVec_2022 <= _zz_regVec_0;
          end
          if(_zz_1[2023]) begin
            regVec_2023 <= _zz_regVec_0;
          end
          if(_zz_1[2024]) begin
            regVec_2024 <= _zz_regVec_0;
          end
          if(_zz_1[2025]) begin
            regVec_2025 <= _zz_regVec_0;
          end
          if(_zz_1[2026]) begin
            regVec_2026 <= _zz_regVec_0;
          end
          if(_zz_1[2027]) begin
            regVec_2027 <= _zz_regVec_0;
          end
          if(_zz_1[2028]) begin
            regVec_2028 <= _zz_regVec_0;
          end
          if(_zz_1[2029]) begin
            regVec_2029 <= _zz_regVec_0;
          end
          if(_zz_1[2030]) begin
            regVec_2030 <= _zz_regVec_0;
          end
          if(_zz_1[2031]) begin
            regVec_2031 <= _zz_regVec_0;
          end
          if(_zz_1[2032]) begin
            regVec_2032 <= _zz_regVec_0;
          end
          if(_zz_1[2033]) begin
            regVec_2033 <= _zz_regVec_0;
          end
          if(_zz_1[2034]) begin
            regVec_2034 <= _zz_regVec_0;
          end
          if(_zz_1[2035]) begin
            regVec_2035 <= _zz_regVec_0;
          end
          if(_zz_1[2036]) begin
            regVec_2036 <= _zz_regVec_0;
          end
          if(_zz_1[2037]) begin
            regVec_2037 <= _zz_regVec_0;
          end
          if(_zz_1[2038]) begin
            regVec_2038 <= _zz_regVec_0;
          end
          if(_zz_1[2039]) begin
            regVec_2039 <= _zz_regVec_0;
          end
          if(_zz_1[2040]) begin
            regVec_2040 <= _zz_regVec_0;
          end
          if(_zz_1[2041]) begin
            regVec_2041 <= _zz_regVec_0;
          end
          if(_zz_1[2042]) begin
            regVec_2042 <= _zz_regVec_0;
          end
          if(_zz_1[2043]) begin
            regVec_2043 <= _zz_regVec_0;
          end
          if(_zz_1[2044]) begin
            regVec_2044 <= _zz_regVec_0;
          end
          if(_zz_1[2045]) begin
            regVec_2045 <= _zz_regVec_0;
          end
          if(_zz_1[2046]) begin
            regVec_2046 <= _zz_regVec_0;
          end
          if(_zz_1[2047]) begin
            regVec_2047 <= _zz_regVec_0;
          end
          if(_zz_1[2048]) begin
            regVec_2048 <= _zz_regVec_0;
          end
          if(_zz_1[2049]) begin
            regVec_2049 <= _zz_regVec_0;
          end
          if(_zz_1[2050]) begin
            regVec_2050 <= _zz_regVec_0;
          end
          if(_zz_1[2051]) begin
            regVec_2051 <= _zz_regVec_0;
          end
          if(_zz_1[2052]) begin
            regVec_2052 <= _zz_regVec_0;
          end
          if(_zz_1[2053]) begin
            regVec_2053 <= _zz_regVec_0;
          end
          if(_zz_1[2054]) begin
            regVec_2054 <= _zz_regVec_0;
          end
          if(_zz_1[2055]) begin
            regVec_2055 <= _zz_regVec_0;
          end
          if(_zz_1[2056]) begin
            regVec_2056 <= _zz_regVec_0;
          end
          if(_zz_1[2057]) begin
            regVec_2057 <= _zz_regVec_0;
          end
          if(_zz_1[2058]) begin
            regVec_2058 <= _zz_regVec_0;
          end
          if(_zz_1[2059]) begin
            regVec_2059 <= _zz_regVec_0;
          end
          if(_zz_1[2060]) begin
            regVec_2060 <= _zz_regVec_0;
          end
          if(_zz_1[2061]) begin
            regVec_2061 <= _zz_regVec_0;
          end
          if(_zz_1[2062]) begin
            regVec_2062 <= _zz_regVec_0;
          end
          if(_zz_1[2063]) begin
            regVec_2063 <= _zz_regVec_0;
          end
          if(_zz_1[2064]) begin
            regVec_2064 <= _zz_regVec_0;
          end
          if(_zz_1[2065]) begin
            regVec_2065 <= _zz_regVec_0;
          end
          if(_zz_1[2066]) begin
            regVec_2066 <= _zz_regVec_0;
          end
          if(_zz_1[2067]) begin
            regVec_2067 <= _zz_regVec_0;
          end
          if(_zz_1[2068]) begin
            regVec_2068 <= _zz_regVec_0;
          end
          if(_zz_1[2069]) begin
            regVec_2069 <= _zz_regVec_0;
          end
          if(_zz_1[2070]) begin
            regVec_2070 <= _zz_regVec_0;
          end
          if(_zz_1[2071]) begin
            regVec_2071 <= _zz_regVec_0;
          end
          if(_zz_1[2072]) begin
            regVec_2072 <= _zz_regVec_0;
          end
          if(_zz_1[2073]) begin
            regVec_2073 <= _zz_regVec_0;
          end
          if(_zz_1[2074]) begin
            regVec_2074 <= _zz_regVec_0;
          end
          if(_zz_1[2075]) begin
            regVec_2075 <= _zz_regVec_0;
          end
          if(_zz_1[2076]) begin
            regVec_2076 <= _zz_regVec_0;
          end
          if(_zz_1[2077]) begin
            regVec_2077 <= _zz_regVec_0;
          end
          if(_zz_1[2078]) begin
            regVec_2078 <= _zz_regVec_0;
          end
          if(_zz_1[2079]) begin
            regVec_2079 <= _zz_regVec_0;
          end
          if(_zz_1[2080]) begin
            regVec_2080 <= _zz_regVec_0;
          end
          if(_zz_1[2081]) begin
            regVec_2081 <= _zz_regVec_0;
          end
          if(_zz_1[2082]) begin
            regVec_2082 <= _zz_regVec_0;
          end
          if(_zz_1[2083]) begin
            regVec_2083 <= _zz_regVec_0;
          end
          if(_zz_1[2084]) begin
            regVec_2084 <= _zz_regVec_0;
          end
          if(_zz_1[2085]) begin
            regVec_2085 <= _zz_regVec_0;
          end
          if(_zz_1[2086]) begin
            regVec_2086 <= _zz_regVec_0;
          end
          if(_zz_1[2087]) begin
            regVec_2087 <= _zz_regVec_0;
          end
          if(_zz_1[2088]) begin
            regVec_2088 <= _zz_regVec_0;
          end
          if(_zz_1[2089]) begin
            regVec_2089 <= _zz_regVec_0;
          end
          if(_zz_1[2090]) begin
            regVec_2090 <= _zz_regVec_0;
          end
          if(_zz_1[2091]) begin
            regVec_2091 <= _zz_regVec_0;
          end
          if(_zz_1[2092]) begin
            regVec_2092 <= _zz_regVec_0;
          end
          if(_zz_1[2093]) begin
            regVec_2093 <= _zz_regVec_0;
          end
          if(_zz_1[2094]) begin
            regVec_2094 <= _zz_regVec_0;
          end
          if(_zz_1[2095]) begin
            regVec_2095 <= _zz_regVec_0;
          end
          if(_zz_1[2096]) begin
            regVec_2096 <= _zz_regVec_0;
          end
          if(_zz_1[2097]) begin
            regVec_2097 <= _zz_regVec_0;
          end
          if(_zz_1[2098]) begin
            regVec_2098 <= _zz_regVec_0;
          end
          if(_zz_1[2099]) begin
            regVec_2099 <= _zz_regVec_0;
          end
          if(_zz_1[2100]) begin
            regVec_2100 <= _zz_regVec_0;
          end
          if(_zz_1[2101]) begin
            regVec_2101 <= _zz_regVec_0;
          end
          if(_zz_1[2102]) begin
            regVec_2102 <= _zz_regVec_0;
          end
          if(_zz_1[2103]) begin
            regVec_2103 <= _zz_regVec_0;
          end
          if(_zz_1[2104]) begin
            regVec_2104 <= _zz_regVec_0;
          end
          if(_zz_1[2105]) begin
            regVec_2105 <= _zz_regVec_0;
          end
          if(_zz_1[2106]) begin
            regVec_2106 <= _zz_regVec_0;
          end
          if(_zz_1[2107]) begin
            regVec_2107 <= _zz_regVec_0;
          end
          if(_zz_1[2108]) begin
            regVec_2108 <= _zz_regVec_0;
          end
          if(_zz_1[2109]) begin
            regVec_2109 <= _zz_regVec_0;
          end
          if(_zz_1[2110]) begin
            regVec_2110 <= _zz_regVec_0;
          end
          if(_zz_1[2111]) begin
            regVec_2111 <= _zz_regVec_0;
          end
          if(_zz_1[2112]) begin
            regVec_2112 <= _zz_regVec_0;
          end
          if(_zz_1[2113]) begin
            regVec_2113 <= _zz_regVec_0;
          end
          if(_zz_1[2114]) begin
            regVec_2114 <= _zz_regVec_0;
          end
          if(_zz_1[2115]) begin
            regVec_2115 <= _zz_regVec_0;
          end
          if(_zz_1[2116]) begin
            regVec_2116 <= _zz_regVec_0;
          end
          if(_zz_1[2117]) begin
            regVec_2117 <= _zz_regVec_0;
          end
          if(_zz_1[2118]) begin
            regVec_2118 <= _zz_regVec_0;
          end
          if(_zz_1[2119]) begin
            regVec_2119 <= _zz_regVec_0;
          end
          if(_zz_1[2120]) begin
            regVec_2120 <= _zz_regVec_0;
          end
          if(_zz_1[2121]) begin
            regVec_2121 <= _zz_regVec_0;
          end
          if(_zz_1[2122]) begin
            regVec_2122 <= _zz_regVec_0;
          end
          if(_zz_1[2123]) begin
            regVec_2123 <= _zz_regVec_0;
          end
          if(_zz_1[2124]) begin
            regVec_2124 <= _zz_regVec_0;
          end
          if(_zz_1[2125]) begin
            regVec_2125 <= _zz_regVec_0;
          end
          if(_zz_1[2126]) begin
            regVec_2126 <= _zz_regVec_0;
          end
          if(_zz_1[2127]) begin
            regVec_2127 <= _zz_regVec_0;
          end
          if(_zz_1[2128]) begin
            regVec_2128 <= _zz_regVec_0;
          end
          if(_zz_1[2129]) begin
            regVec_2129 <= _zz_regVec_0;
          end
          if(_zz_1[2130]) begin
            regVec_2130 <= _zz_regVec_0;
          end
          if(_zz_1[2131]) begin
            regVec_2131 <= _zz_regVec_0;
          end
          if(_zz_1[2132]) begin
            regVec_2132 <= _zz_regVec_0;
          end
          if(_zz_1[2133]) begin
            regVec_2133 <= _zz_regVec_0;
          end
          if(_zz_1[2134]) begin
            regVec_2134 <= _zz_regVec_0;
          end
          if(_zz_1[2135]) begin
            regVec_2135 <= _zz_regVec_0;
          end
          if(_zz_1[2136]) begin
            regVec_2136 <= _zz_regVec_0;
          end
          if(_zz_1[2137]) begin
            regVec_2137 <= _zz_regVec_0;
          end
          if(_zz_1[2138]) begin
            regVec_2138 <= _zz_regVec_0;
          end
          if(_zz_1[2139]) begin
            regVec_2139 <= _zz_regVec_0;
          end
          if(_zz_1[2140]) begin
            regVec_2140 <= _zz_regVec_0;
          end
          if(_zz_1[2141]) begin
            regVec_2141 <= _zz_regVec_0;
          end
          if(_zz_1[2142]) begin
            regVec_2142 <= _zz_regVec_0;
          end
          if(_zz_1[2143]) begin
            regVec_2143 <= _zz_regVec_0;
          end
          if(_zz_1[2144]) begin
            regVec_2144 <= _zz_regVec_0;
          end
          if(_zz_1[2145]) begin
            regVec_2145 <= _zz_regVec_0;
          end
          if(_zz_1[2146]) begin
            regVec_2146 <= _zz_regVec_0;
          end
          if(_zz_1[2147]) begin
            regVec_2147 <= _zz_regVec_0;
          end
          if(_zz_1[2148]) begin
            regVec_2148 <= _zz_regVec_0;
          end
          if(_zz_1[2149]) begin
            regVec_2149 <= _zz_regVec_0;
          end
          if(_zz_1[2150]) begin
            regVec_2150 <= _zz_regVec_0;
          end
          if(_zz_1[2151]) begin
            regVec_2151 <= _zz_regVec_0;
          end
          if(_zz_1[2152]) begin
            regVec_2152 <= _zz_regVec_0;
          end
          if(_zz_1[2153]) begin
            regVec_2153 <= _zz_regVec_0;
          end
          if(_zz_1[2154]) begin
            regVec_2154 <= _zz_regVec_0;
          end
          if(_zz_1[2155]) begin
            regVec_2155 <= _zz_regVec_0;
          end
          if(_zz_1[2156]) begin
            regVec_2156 <= _zz_regVec_0;
          end
          if(_zz_1[2157]) begin
            regVec_2157 <= _zz_regVec_0;
          end
          if(_zz_1[2158]) begin
            regVec_2158 <= _zz_regVec_0;
          end
          if(_zz_1[2159]) begin
            regVec_2159 <= _zz_regVec_0;
          end
          if(_zz_1[2160]) begin
            regVec_2160 <= _zz_regVec_0;
          end
          if(_zz_1[2161]) begin
            regVec_2161 <= _zz_regVec_0;
          end
          if(_zz_1[2162]) begin
            regVec_2162 <= _zz_regVec_0;
          end
          if(_zz_1[2163]) begin
            regVec_2163 <= _zz_regVec_0;
          end
          if(_zz_1[2164]) begin
            regVec_2164 <= _zz_regVec_0;
          end
          if(_zz_1[2165]) begin
            regVec_2165 <= _zz_regVec_0;
          end
          if(_zz_1[2166]) begin
            regVec_2166 <= _zz_regVec_0;
          end
          if(_zz_1[2167]) begin
            regVec_2167 <= _zz_regVec_0;
          end
          if(_zz_1[2168]) begin
            regVec_2168 <= _zz_regVec_0;
          end
          if(_zz_1[2169]) begin
            regVec_2169 <= _zz_regVec_0;
          end
          if(_zz_1[2170]) begin
            regVec_2170 <= _zz_regVec_0;
          end
          if(_zz_1[2171]) begin
            regVec_2171 <= _zz_regVec_0;
          end
          if(_zz_1[2172]) begin
            regVec_2172 <= _zz_regVec_0;
          end
          if(_zz_1[2173]) begin
            regVec_2173 <= _zz_regVec_0;
          end
          if(_zz_1[2174]) begin
            regVec_2174 <= _zz_regVec_0;
          end
          if(_zz_1[2175]) begin
            regVec_2175 <= _zz_regVec_0;
          end
          if(_zz_1[2176]) begin
            regVec_2176 <= _zz_regVec_0;
          end
          if(_zz_1[2177]) begin
            regVec_2177 <= _zz_regVec_0;
          end
          if(_zz_1[2178]) begin
            regVec_2178 <= _zz_regVec_0;
          end
          if(_zz_1[2179]) begin
            regVec_2179 <= _zz_regVec_0;
          end
          if(_zz_1[2180]) begin
            regVec_2180 <= _zz_regVec_0;
          end
          if(_zz_1[2181]) begin
            regVec_2181 <= _zz_regVec_0;
          end
          if(_zz_1[2182]) begin
            regVec_2182 <= _zz_regVec_0;
          end
          if(_zz_1[2183]) begin
            regVec_2183 <= _zz_regVec_0;
          end
          if(_zz_1[2184]) begin
            regVec_2184 <= _zz_regVec_0;
          end
          if(_zz_1[2185]) begin
            regVec_2185 <= _zz_regVec_0;
          end
          if(_zz_1[2186]) begin
            regVec_2186 <= _zz_regVec_0;
          end
          if(_zz_1[2187]) begin
            regVec_2187 <= _zz_regVec_0;
          end
          if(_zz_1[2188]) begin
            regVec_2188 <= _zz_regVec_0;
          end
          if(_zz_1[2189]) begin
            regVec_2189 <= _zz_regVec_0;
          end
          if(_zz_1[2190]) begin
            regVec_2190 <= _zz_regVec_0;
          end
          if(_zz_1[2191]) begin
            regVec_2191 <= _zz_regVec_0;
          end
          if(_zz_1[2192]) begin
            regVec_2192 <= _zz_regVec_0;
          end
          if(_zz_1[2193]) begin
            regVec_2193 <= _zz_regVec_0;
          end
          if(_zz_1[2194]) begin
            regVec_2194 <= _zz_regVec_0;
          end
          if(_zz_1[2195]) begin
            regVec_2195 <= _zz_regVec_0;
          end
          if(_zz_1[2196]) begin
            regVec_2196 <= _zz_regVec_0;
          end
          if(_zz_1[2197]) begin
            regVec_2197 <= _zz_regVec_0;
          end
          if(_zz_1[2198]) begin
            regVec_2198 <= _zz_regVec_0;
          end
          if(_zz_1[2199]) begin
            regVec_2199 <= _zz_regVec_0;
          end
          if(_zz_1[2200]) begin
            regVec_2200 <= _zz_regVec_0;
          end
          if(_zz_1[2201]) begin
            regVec_2201 <= _zz_regVec_0;
          end
          if(_zz_1[2202]) begin
            regVec_2202 <= _zz_regVec_0;
          end
          if(_zz_1[2203]) begin
            regVec_2203 <= _zz_regVec_0;
          end
          if(_zz_1[2204]) begin
            regVec_2204 <= _zz_regVec_0;
          end
          if(_zz_1[2205]) begin
            regVec_2205 <= _zz_regVec_0;
          end
          if(_zz_1[2206]) begin
            regVec_2206 <= _zz_regVec_0;
          end
          if(_zz_1[2207]) begin
            regVec_2207 <= _zz_regVec_0;
          end
          if(_zz_1[2208]) begin
            regVec_2208 <= _zz_regVec_0;
          end
          if(_zz_1[2209]) begin
            regVec_2209 <= _zz_regVec_0;
          end
          if(_zz_1[2210]) begin
            regVec_2210 <= _zz_regVec_0;
          end
          if(_zz_1[2211]) begin
            regVec_2211 <= _zz_regVec_0;
          end
          if(_zz_1[2212]) begin
            regVec_2212 <= _zz_regVec_0;
          end
          if(_zz_1[2213]) begin
            regVec_2213 <= _zz_regVec_0;
          end
          if(_zz_1[2214]) begin
            regVec_2214 <= _zz_regVec_0;
          end
          if(_zz_1[2215]) begin
            regVec_2215 <= _zz_regVec_0;
          end
          if(_zz_1[2216]) begin
            regVec_2216 <= _zz_regVec_0;
          end
          if(_zz_1[2217]) begin
            regVec_2217 <= _zz_regVec_0;
          end
          if(_zz_1[2218]) begin
            regVec_2218 <= _zz_regVec_0;
          end
          if(_zz_1[2219]) begin
            regVec_2219 <= _zz_regVec_0;
          end
          if(_zz_1[2220]) begin
            regVec_2220 <= _zz_regVec_0;
          end
          if(_zz_1[2221]) begin
            regVec_2221 <= _zz_regVec_0;
          end
          if(_zz_1[2222]) begin
            regVec_2222 <= _zz_regVec_0;
          end
          if(_zz_1[2223]) begin
            regVec_2223 <= _zz_regVec_0;
          end
          if(_zz_1[2224]) begin
            regVec_2224 <= _zz_regVec_0;
          end
          if(_zz_1[2225]) begin
            regVec_2225 <= _zz_regVec_0;
          end
          if(_zz_1[2226]) begin
            regVec_2226 <= _zz_regVec_0;
          end
          if(_zz_1[2227]) begin
            regVec_2227 <= _zz_regVec_0;
          end
          if(_zz_1[2228]) begin
            regVec_2228 <= _zz_regVec_0;
          end
          if(_zz_1[2229]) begin
            regVec_2229 <= _zz_regVec_0;
          end
          if(_zz_1[2230]) begin
            regVec_2230 <= _zz_regVec_0;
          end
          if(_zz_1[2231]) begin
            regVec_2231 <= _zz_regVec_0;
          end
          if(_zz_1[2232]) begin
            regVec_2232 <= _zz_regVec_0;
          end
          if(_zz_1[2233]) begin
            regVec_2233 <= _zz_regVec_0;
          end
          if(_zz_1[2234]) begin
            regVec_2234 <= _zz_regVec_0;
          end
          if(_zz_1[2235]) begin
            regVec_2235 <= _zz_regVec_0;
          end
          if(_zz_1[2236]) begin
            regVec_2236 <= _zz_regVec_0;
          end
          if(_zz_1[2237]) begin
            regVec_2237 <= _zz_regVec_0;
          end
          if(_zz_1[2238]) begin
            regVec_2238 <= _zz_regVec_0;
          end
          if(_zz_1[2239]) begin
            regVec_2239 <= _zz_regVec_0;
          end
          if(_zz_1[2240]) begin
            regVec_2240 <= _zz_regVec_0;
          end
          if(_zz_1[2241]) begin
            regVec_2241 <= _zz_regVec_0;
          end
          if(_zz_1[2242]) begin
            regVec_2242 <= _zz_regVec_0;
          end
          if(_zz_1[2243]) begin
            regVec_2243 <= _zz_regVec_0;
          end
          if(_zz_1[2244]) begin
            regVec_2244 <= _zz_regVec_0;
          end
          if(_zz_1[2245]) begin
            regVec_2245 <= _zz_regVec_0;
          end
          if(_zz_1[2246]) begin
            regVec_2246 <= _zz_regVec_0;
          end
          if(_zz_1[2247]) begin
            regVec_2247 <= _zz_regVec_0;
          end
          if(_zz_1[2248]) begin
            regVec_2248 <= _zz_regVec_0;
          end
          if(_zz_1[2249]) begin
            regVec_2249 <= _zz_regVec_0;
          end
          if(_zz_1[2250]) begin
            regVec_2250 <= _zz_regVec_0;
          end
          if(_zz_1[2251]) begin
            regVec_2251 <= _zz_regVec_0;
          end
          if(_zz_1[2252]) begin
            regVec_2252 <= _zz_regVec_0;
          end
          if(_zz_1[2253]) begin
            regVec_2253 <= _zz_regVec_0;
          end
          if(_zz_1[2254]) begin
            regVec_2254 <= _zz_regVec_0;
          end
          if(_zz_1[2255]) begin
            regVec_2255 <= _zz_regVec_0;
          end
          if(_zz_1[2256]) begin
            regVec_2256 <= _zz_regVec_0;
          end
          if(_zz_1[2257]) begin
            regVec_2257 <= _zz_regVec_0;
          end
          if(_zz_1[2258]) begin
            regVec_2258 <= _zz_regVec_0;
          end
          if(_zz_1[2259]) begin
            regVec_2259 <= _zz_regVec_0;
          end
          if(_zz_1[2260]) begin
            regVec_2260 <= _zz_regVec_0;
          end
          if(_zz_1[2261]) begin
            regVec_2261 <= _zz_regVec_0;
          end
          if(_zz_1[2262]) begin
            regVec_2262 <= _zz_regVec_0;
          end
          if(_zz_1[2263]) begin
            regVec_2263 <= _zz_regVec_0;
          end
          if(_zz_1[2264]) begin
            regVec_2264 <= _zz_regVec_0;
          end
          if(_zz_1[2265]) begin
            regVec_2265 <= _zz_regVec_0;
          end
          if(_zz_1[2266]) begin
            regVec_2266 <= _zz_regVec_0;
          end
          if(_zz_1[2267]) begin
            regVec_2267 <= _zz_regVec_0;
          end
          if(_zz_1[2268]) begin
            regVec_2268 <= _zz_regVec_0;
          end
          if(_zz_1[2269]) begin
            regVec_2269 <= _zz_regVec_0;
          end
          if(_zz_1[2270]) begin
            regVec_2270 <= _zz_regVec_0;
          end
          if(_zz_1[2271]) begin
            regVec_2271 <= _zz_regVec_0;
          end
          if(_zz_1[2272]) begin
            regVec_2272 <= _zz_regVec_0;
          end
          if(_zz_1[2273]) begin
            regVec_2273 <= _zz_regVec_0;
          end
          if(_zz_1[2274]) begin
            regVec_2274 <= _zz_regVec_0;
          end
          if(_zz_1[2275]) begin
            regVec_2275 <= _zz_regVec_0;
          end
          if(_zz_1[2276]) begin
            regVec_2276 <= _zz_regVec_0;
          end
          if(_zz_1[2277]) begin
            regVec_2277 <= _zz_regVec_0;
          end
          if(_zz_1[2278]) begin
            regVec_2278 <= _zz_regVec_0;
          end
          if(_zz_1[2279]) begin
            regVec_2279 <= _zz_regVec_0;
          end
          if(_zz_1[2280]) begin
            regVec_2280 <= _zz_regVec_0;
          end
          if(_zz_1[2281]) begin
            regVec_2281 <= _zz_regVec_0;
          end
          if(_zz_1[2282]) begin
            regVec_2282 <= _zz_regVec_0;
          end
          if(_zz_1[2283]) begin
            regVec_2283 <= _zz_regVec_0;
          end
          if(_zz_1[2284]) begin
            regVec_2284 <= _zz_regVec_0;
          end
          if(_zz_1[2285]) begin
            regVec_2285 <= _zz_regVec_0;
          end
          if(_zz_1[2286]) begin
            regVec_2286 <= _zz_regVec_0;
          end
          if(_zz_1[2287]) begin
            regVec_2287 <= _zz_regVec_0;
          end
          if(_zz_1[2288]) begin
            regVec_2288 <= _zz_regVec_0;
          end
          if(_zz_1[2289]) begin
            regVec_2289 <= _zz_regVec_0;
          end
          if(_zz_1[2290]) begin
            regVec_2290 <= _zz_regVec_0;
          end
          if(_zz_1[2291]) begin
            regVec_2291 <= _zz_regVec_0;
          end
          if(_zz_1[2292]) begin
            regVec_2292 <= _zz_regVec_0;
          end
          if(_zz_1[2293]) begin
            regVec_2293 <= _zz_regVec_0;
          end
          if(_zz_1[2294]) begin
            regVec_2294 <= _zz_regVec_0;
          end
          if(_zz_1[2295]) begin
            regVec_2295 <= _zz_regVec_0;
          end
          if(_zz_1[2296]) begin
            regVec_2296 <= _zz_regVec_0;
          end
          if(_zz_1[2297]) begin
            regVec_2297 <= _zz_regVec_0;
          end
          if(_zz_1[2298]) begin
            regVec_2298 <= _zz_regVec_0;
          end
          if(_zz_1[2299]) begin
            regVec_2299 <= _zz_regVec_0;
          end
          if(_zz_1[2300]) begin
            regVec_2300 <= _zz_regVec_0;
          end
          if(_zz_1[2301]) begin
            regVec_2301 <= _zz_regVec_0;
          end
          if(_zz_1[2302]) begin
            regVec_2302 <= _zz_regVec_0;
          end
          if(_zz_1[2303]) begin
            regVec_2303 <= _zz_regVec_0;
          end
          if(_zz_1[2304]) begin
            regVec_2304 <= _zz_regVec_0;
          end
          if(_zz_1[2305]) begin
            regVec_2305 <= _zz_regVec_0;
          end
          if(_zz_1[2306]) begin
            regVec_2306 <= _zz_regVec_0;
          end
          if(_zz_1[2307]) begin
            regVec_2307 <= _zz_regVec_0;
          end
          if(_zz_1[2308]) begin
            regVec_2308 <= _zz_regVec_0;
          end
          if(_zz_1[2309]) begin
            regVec_2309 <= _zz_regVec_0;
          end
          if(_zz_1[2310]) begin
            regVec_2310 <= _zz_regVec_0;
          end
          if(_zz_1[2311]) begin
            regVec_2311 <= _zz_regVec_0;
          end
          if(_zz_1[2312]) begin
            regVec_2312 <= _zz_regVec_0;
          end
          if(_zz_1[2313]) begin
            regVec_2313 <= _zz_regVec_0;
          end
          if(_zz_1[2314]) begin
            regVec_2314 <= _zz_regVec_0;
          end
          if(_zz_1[2315]) begin
            regVec_2315 <= _zz_regVec_0;
          end
          if(_zz_1[2316]) begin
            regVec_2316 <= _zz_regVec_0;
          end
          if(_zz_1[2317]) begin
            regVec_2317 <= _zz_regVec_0;
          end
          if(_zz_1[2318]) begin
            regVec_2318 <= _zz_regVec_0;
          end
          if(_zz_1[2319]) begin
            regVec_2319 <= _zz_regVec_0;
          end
          if(_zz_1[2320]) begin
            regVec_2320 <= _zz_regVec_0;
          end
          if(_zz_1[2321]) begin
            regVec_2321 <= _zz_regVec_0;
          end
          if(_zz_1[2322]) begin
            regVec_2322 <= _zz_regVec_0;
          end
          if(_zz_1[2323]) begin
            regVec_2323 <= _zz_regVec_0;
          end
          if(_zz_1[2324]) begin
            regVec_2324 <= _zz_regVec_0;
          end
          if(_zz_1[2325]) begin
            regVec_2325 <= _zz_regVec_0;
          end
          if(_zz_1[2326]) begin
            regVec_2326 <= _zz_regVec_0;
          end
          if(_zz_1[2327]) begin
            regVec_2327 <= _zz_regVec_0;
          end
          if(_zz_1[2328]) begin
            regVec_2328 <= _zz_regVec_0;
          end
          if(_zz_1[2329]) begin
            regVec_2329 <= _zz_regVec_0;
          end
          if(_zz_1[2330]) begin
            regVec_2330 <= _zz_regVec_0;
          end
          if(_zz_1[2331]) begin
            regVec_2331 <= _zz_regVec_0;
          end
          if(_zz_1[2332]) begin
            regVec_2332 <= _zz_regVec_0;
          end
          if(_zz_1[2333]) begin
            regVec_2333 <= _zz_regVec_0;
          end
          if(_zz_1[2334]) begin
            regVec_2334 <= _zz_regVec_0;
          end
          if(_zz_1[2335]) begin
            regVec_2335 <= _zz_regVec_0;
          end
          if(_zz_1[2336]) begin
            regVec_2336 <= _zz_regVec_0;
          end
          if(_zz_1[2337]) begin
            regVec_2337 <= _zz_regVec_0;
          end
          if(_zz_1[2338]) begin
            regVec_2338 <= _zz_regVec_0;
          end
          if(_zz_1[2339]) begin
            regVec_2339 <= _zz_regVec_0;
          end
          if(_zz_1[2340]) begin
            regVec_2340 <= _zz_regVec_0;
          end
          if(_zz_1[2341]) begin
            regVec_2341 <= _zz_regVec_0;
          end
          if(_zz_1[2342]) begin
            regVec_2342 <= _zz_regVec_0;
          end
          if(_zz_1[2343]) begin
            regVec_2343 <= _zz_regVec_0;
          end
          if(_zz_1[2344]) begin
            regVec_2344 <= _zz_regVec_0;
          end
          if(_zz_1[2345]) begin
            regVec_2345 <= _zz_regVec_0;
          end
          if(_zz_1[2346]) begin
            regVec_2346 <= _zz_regVec_0;
          end
          if(_zz_1[2347]) begin
            regVec_2347 <= _zz_regVec_0;
          end
          if(_zz_1[2348]) begin
            regVec_2348 <= _zz_regVec_0;
          end
          if(_zz_1[2349]) begin
            regVec_2349 <= _zz_regVec_0;
          end
          if(_zz_1[2350]) begin
            regVec_2350 <= _zz_regVec_0;
          end
          if(_zz_1[2351]) begin
            regVec_2351 <= _zz_regVec_0;
          end
          if(_zz_1[2352]) begin
            regVec_2352 <= _zz_regVec_0;
          end
          if(_zz_1[2353]) begin
            regVec_2353 <= _zz_regVec_0;
          end
          if(_zz_1[2354]) begin
            regVec_2354 <= _zz_regVec_0;
          end
          if(_zz_1[2355]) begin
            regVec_2355 <= _zz_regVec_0;
          end
          if(_zz_1[2356]) begin
            regVec_2356 <= _zz_regVec_0;
          end
          if(_zz_1[2357]) begin
            regVec_2357 <= _zz_regVec_0;
          end
          if(_zz_1[2358]) begin
            regVec_2358 <= _zz_regVec_0;
          end
          if(_zz_1[2359]) begin
            regVec_2359 <= _zz_regVec_0;
          end
          if(_zz_1[2360]) begin
            regVec_2360 <= _zz_regVec_0;
          end
          if(_zz_1[2361]) begin
            regVec_2361 <= _zz_regVec_0;
          end
          if(_zz_1[2362]) begin
            regVec_2362 <= _zz_regVec_0;
          end
          if(_zz_1[2363]) begin
            regVec_2363 <= _zz_regVec_0;
          end
          if(_zz_1[2364]) begin
            regVec_2364 <= _zz_regVec_0;
          end
          if(_zz_1[2365]) begin
            regVec_2365 <= _zz_regVec_0;
          end
          if(_zz_1[2366]) begin
            regVec_2366 <= _zz_regVec_0;
          end
          if(_zz_1[2367]) begin
            regVec_2367 <= _zz_regVec_0;
          end
          if(_zz_1[2368]) begin
            regVec_2368 <= _zz_regVec_0;
          end
          if(_zz_1[2369]) begin
            regVec_2369 <= _zz_regVec_0;
          end
          if(_zz_1[2370]) begin
            regVec_2370 <= _zz_regVec_0;
          end
          if(_zz_1[2371]) begin
            regVec_2371 <= _zz_regVec_0;
          end
          if(_zz_1[2372]) begin
            regVec_2372 <= _zz_regVec_0;
          end
          if(_zz_1[2373]) begin
            regVec_2373 <= _zz_regVec_0;
          end
          if(_zz_1[2374]) begin
            regVec_2374 <= _zz_regVec_0;
          end
          if(_zz_1[2375]) begin
            regVec_2375 <= _zz_regVec_0;
          end
          if(_zz_1[2376]) begin
            regVec_2376 <= _zz_regVec_0;
          end
          if(_zz_1[2377]) begin
            regVec_2377 <= _zz_regVec_0;
          end
          if(_zz_1[2378]) begin
            regVec_2378 <= _zz_regVec_0;
          end
          if(_zz_1[2379]) begin
            regVec_2379 <= _zz_regVec_0;
          end
          if(_zz_1[2380]) begin
            regVec_2380 <= _zz_regVec_0;
          end
          if(_zz_1[2381]) begin
            regVec_2381 <= _zz_regVec_0;
          end
          if(_zz_1[2382]) begin
            regVec_2382 <= _zz_regVec_0;
          end
          if(_zz_1[2383]) begin
            regVec_2383 <= _zz_regVec_0;
          end
          if(_zz_1[2384]) begin
            regVec_2384 <= _zz_regVec_0;
          end
          if(_zz_1[2385]) begin
            regVec_2385 <= _zz_regVec_0;
          end
          if(_zz_1[2386]) begin
            regVec_2386 <= _zz_regVec_0;
          end
          if(_zz_1[2387]) begin
            regVec_2387 <= _zz_regVec_0;
          end
          if(_zz_1[2388]) begin
            regVec_2388 <= _zz_regVec_0;
          end
          if(_zz_1[2389]) begin
            regVec_2389 <= _zz_regVec_0;
          end
          if(_zz_1[2390]) begin
            regVec_2390 <= _zz_regVec_0;
          end
          if(_zz_1[2391]) begin
            regVec_2391 <= _zz_regVec_0;
          end
          if(_zz_1[2392]) begin
            regVec_2392 <= _zz_regVec_0;
          end
          if(_zz_1[2393]) begin
            regVec_2393 <= _zz_regVec_0;
          end
          if(_zz_1[2394]) begin
            regVec_2394 <= _zz_regVec_0;
          end
          if(_zz_1[2395]) begin
            regVec_2395 <= _zz_regVec_0;
          end
          if(_zz_1[2396]) begin
            regVec_2396 <= _zz_regVec_0;
          end
          if(_zz_1[2397]) begin
            regVec_2397 <= _zz_regVec_0;
          end
          if(_zz_1[2398]) begin
            regVec_2398 <= _zz_regVec_0;
          end
          if(_zz_1[2399]) begin
            regVec_2399 <= _zz_regVec_0;
          end
          if(_zz_1[2400]) begin
            regVec_2400 <= _zz_regVec_0;
          end
          if(_zz_1[2401]) begin
            regVec_2401 <= _zz_regVec_0;
          end
          if(_zz_1[2402]) begin
            regVec_2402 <= _zz_regVec_0;
          end
          if(_zz_1[2403]) begin
            regVec_2403 <= _zz_regVec_0;
          end
          if(_zz_1[2404]) begin
            regVec_2404 <= _zz_regVec_0;
          end
          if(_zz_1[2405]) begin
            regVec_2405 <= _zz_regVec_0;
          end
          if(_zz_1[2406]) begin
            regVec_2406 <= _zz_regVec_0;
          end
          if(_zz_1[2407]) begin
            regVec_2407 <= _zz_regVec_0;
          end
          if(_zz_1[2408]) begin
            regVec_2408 <= _zz_regVec_0;
          end
          if(_zz_1[2409]) begin
            regVec_2409 <= _zz_regVec_0;
          end
          if(_zz_1[2410]) begin
            regVec_2410 <= _zz_regVec_0;
          end
          if(_zz_1[2411]) begin
            regVec_2411 <= _zz_regVec_0;
          end
          if(_zz_1[2412]) begin
            regVec_2412 <= _zz_regVec_0;
          end
          if(_zz_1[2413]) begin
            regVec_2413 <= _zz_regVec_0;
          end
          if(_zz_1[2414]) begin
            regVec_2414 <= _zz_regVec_0;
          end
          if(_zz_1[2415]) begin
            regVec_2415 <= _zz_regVec_0;
          end
          if(_zz_1[2416]) begin
            regVec_2416 <= _zz_regVec_0;
          end
          if(_zz_1[2417]) begin
            regVec_2417 <= _zz_regVec_0;
          end
          if(_zz_1[2418]) begin
            regVec_2418 <= _zz_regVec_0;
          end
          if(_zz_1[2419]) begin
            regVec_2419 <= _zz_regVec_0;
          end
          if(_zz_1[2420]) begin
            regVec_2420 <= _zz_regVec_0;
          end
          if(_zz_1[2421]) begin
            regVec_2421 <= _zz_regVec_0;
          end
          if(_zz_1[2422]) begin
            regVec_2422 <= _zz_regVec_0;
          end
          if(_zz_1[2423]) begin
            regVec_2423 <= _zz_regVec_0;
          end
          if(_zz_1[2424]) begin
            regVec_2424 <= _zz_regVec_0;
          end
          if(_zz_1[2425]) begin
            regVec_2425 <= _zz_regVec_0;
          end
          if(_zz_1[2426]) begin
            regVec_2426 <= _zz_regVec_0;
          end
          if(_zz_1[2427]) begin
            regVec_2427 <= _zz_regVec_0;
          end
          if(_zz_1[2428]) begin
            regVec_2428 <= _zz_regVec_0;
          end
          if(_zz_1[2429]) begin
            regVec_2429 <= _zz_regVec_0;
          end
          if(_zz_1[2430]) begin
            regVec_2430 <= _zz_regVec_0;
          end
          if(_zz_1[2431]) begin
            regVec_2431 <= _zz_regVec_0;
          end
          if(_zz_1[2432]) begin
            regVec_2432 <= _zz_regVec_0;
          end
          if(_zz_1[2433]) begin
            regVec_2433 <= _zz_regVec_0;
          end
          if(_zz_1[2434]) begin
            regVec_2434 <= _zz_regVec_0;
          end
          if(_zz_1[2435]) begin
            regVec_2435 <= _zz_regVec_0;
          end
          if(_zz_1[2436]) begin
            regVec_2436 <= _zz_regVec_0;
          end
          if(_zz_1[2437]) begin
            regVec_2437 <= _zz_regVec_0;
          end
          if(_zz_1[2438]) begin
            regVec_2438 <= _zz_regVec_0;
          end
          if(_zz_1[2439]) begin
            regVec_2439 <= _zz_regVec_0;
          end
          if(_zz_1[2440]) begin
            regVec_2440 <= _zz_regVec_0;
          end
          if(_zz_1[2441]) begin
            regVec_2441 <= _zz_regVec_0;
          end
          if(_zz_1[2442]) begin
            regVec_2442 <= _zz_regVec_0;
          end
          if(_zz_1[2443]) begin
            regVec_2443 <= _zz_regVec_0;
          end
          if(_zz_1[2444]) begin
            regVec_2444 <= _zz_regVec_0;
          end
          if(_zz_1[2445]) begin
            regVec_2445 <= _zz_regVec_0;
          end
          if(_zz_1[2446]) begin
            regVec_2446 <= _zz_regVec_0;
          end
          if(_zz_1[2447]) begin
            regVec_2447 <= _zz_regVec_0;
          end
          if(_zz_1[2448]) begin
            regVec_2448 <= _zz_regVec_0;
          end
          if(_zz_1[2449]) begin
            regVec_2449 <= _zz_regVec_0;
          end
          if(_zz_1[2450]) begin
            regVec_2450 <= _zz_regVec_0;
          end
          if(_zz_1[2451]) begin
            regVec_2451 <= _zz_regVec_0;
          end
          if(_zz_1[2452]) begin
            regVec_2452 <= _zz_regVec_0;
          end
          if(_zz_1[2453]) begin
            regVec_2453 <= _zz_regVec_0;
          end
          if(_zz_1[2454]) begin
            regVec_2454 <= _zz_regVec_0;
          end
          if(_zz_1[2455]) begin
            regVec_2455 <= _zz_regVec_0;
          end
          if(_zz_1[2456]) begin
            regVec_2456 <= _zz_regVec_0;
          end
          if(_zz_1[2457]) begin
            regVec_2457 <= _zz_regVec_0;
          end
          if(_zz_1[2458]) begin
            regVec_2458 <= _zz_regVec_0;
          end
          if(_zz_1[2459]) begin
            regVec_2459 <= _zz_regVec_0;
          end
          if(_zz_1[2460]) begin
            regVec_2460 <= _zz_regVec_0;
          end
          if(_zz_1[2461]) begin
            regVec_2461 <= _zz_regVec_0;
          end
          if(_zz_1[2462]) begin
            regVec_2462 <= _zz_regVec_0;
          end
          if(_zz_1[2463]) begin
            regVec_2463 <= _zz_regVec_0;
          end
          if(_zz_1[2464]) begin
            regVec_2464 <= _zz_regVec_0;
          end
          if(_zz_1[2465]) begin
            regVec_2465 <= _zz_regVec_0;
          end
          if(_zz_1[2466]) begin
            regVec_2466 <= _zz_regVec_0;
          end
          if(_zz_1[2467]) begin
            regVec_2467 <= _zz_regVec_0;
          end
          if(_zz_1[2468]) begin
            regVec_2468 <= _zz_regVec_0;
          end
          if(_zz_1[2469]) begin
            regVec_2469 <= _zz_regVec_0;
          end
          if(_zz_1[2470]) begin
            regVec_2470 <= _zz_regVec_0;
          end
          if(_zz_1[2471]) begin
            regVec_2471 <= _zz_regVec_0;
          end
          if(_zz_1[2472]) begin
            regVec_2472 <= _zz_regVec_0;
          end
          if(_zz_1[2473]) begin
            regVec_2473 <= _zz_regVec_0;
          end
          if(_zz_1[2474]) begin
            regVec_2474 <= _zz_regVec_0;
          end
          if(_zz_1[2475]) begin
            regVec_2475 <= _zz_regVec_0;
          end
          if(_zz_1[2476]) begin
            regVec_2476 <= _zz_regVec_0;
          end
          if(_zz_1[2477]) begin
            regVec_2477 <= _zz_regVec_0;
          end
          if(_zz_1[2478]) begin
            regVec_2478 <= _zz_regVec_0;
          end
          if(_zz_1[2479]) begin
            regVec_2479 <= _zz_regVec_0;
          end
          if(_zz_1[2480]) begin
            regVec_2480 <= _zz_regVec_0;
          end
          if(_zz_1[2481]) begin
            regVec_2481 <= _zz_regVec_0;
          end
          if(_zz_1[2482]) begin
            regVec_2482 <= _zz_regVec_0;
          end
          if(_zz_1[2483]) begin
            regVec_2483 <= _zz_regVec_0;
          end
          if(_zz_1[2484]) begin
            regVec_2484 <= _zz_regVec_0;
          end
          if(_zz_1[2485]) begin
            regVec_2485 <= _zz_regVec_0;
          end
          if(_zz_1[2486]) begin
            regVec_2486 <= _zz_regVec_0;
          end
          if(_zz_1[2487]) begin
            regVec_2487 <= _zz_regVec_0;
          end
          if(_zz_1[2488]) begin
            regVec_2488 <= _zz_regVec_0;
          end
          if(_zz_1[2489]) begin
            regVec_2489 <= _zz_regVec_0;
          end
          if(_zz_1[2490]) begin
            regVec_2490 <= _zz_regVec_0;
          end
          if(_zz_1[2491]) begin
            regVec_2491 <= _zz_regVec_0;
          end
          if(_zz_1[2492]) begin
            regVec_2492 <= _zz_regVec_0;
          end
          if(_zz_1[2493]) begin
            regVec_2493 <= _zz_regVec_0;
          end
          if(_zz_1[2494]) begin
            regVec_2494 <= _zz_regVec_0;
          end
          if(_zz_1[2495]) begin
            regVec_2495 <= _zz_regVec_0;
          end
          if(_zz_1[2496]) begin
            regVec_2496 <= _zz_regVec_0;
          end
          if(_zz_1[2497]) begin
            regVec_2497 <= _zz_regVec_0;
          end
          if(_zz_1[2498]) begin
            regVec_2498 <= _zz_regVec_0;
          end
          if(_zz_1[2499]) begin
            regVec_2499 <= _zz_regVec_0;
          end
          if(_zz_1[2500]) begin
            regVec_2500 <= _zz_regVec_0;
          end
          if(_zz_1[2501]) begin
            regVec_2501 <= _zz_regVec_0;
          end
          if(_zz_1[2502]) begin
            regVec_2502 <= _zz_regVec_0;
          end
          if(_zz_1[2503]) begin
            regVec_2503 <= _zz_regVec_0;
          end
          if(_zz_1[2504]) begin
            regVec_2504 <= _zz_regVec_0;
          end
          if(_zz_1[2505]) begin
            regVec_2505 <= _zz_regVec_0;
          end
          if(_zz_1[2506]) begin
            regVec_2506 <= _zz_regVec_0;
          end
          if(_zz_1[2507]) begin
            regVec_2507 <= _zz_regVec_0;
          end
          if(_zz_1[2508]) begin
            regVec_2508 <= _zz_regVec_0;
          end
          if(_zz_1[2509]) begin
            regVec_2509 <= _zz_regVec_0;
          end
          if(_zz_1[2510]) begin
            regVec_2510 <= _zz_regVec_0;
          end
          if(_zz_1[2511]) begin
            regVec_2511 <= _zz_regVec_0;
          end
          if(_zz_1[2512]) begin
            regVec_2512 <= _zz_regVec_0;
          end
          if(_zz_1[2513]) begin
            regVec_2513 <= _zz_regVec_0;
          end
          if(_zz_1[2514]) begin
            regVec_2514 <= _zz_regVec_0;
          end
          if(_zz_1[2515]) begin
            regVec_2515 <= _zz_regVec_0;
          end
          if(_zz_1[2516]) begin
            regVec_2516 <= _zz_regVec_0;
          end
          if(_zz_1[2517]) begin
            regVec_2517 <= _zz_regVec_0;
          end
          if(_zz_1[2518]) begin
            regVec_2518 <= _zz_regVec_0;
          end
          if(_zz_1[2519]) begin
            regVec_2519 <= _zz_regVec_0;
          end
          if(_zz_1[2520]) begin
            regVec_2520 <= _zz_regVec_0;
          end
          if(_zz_1[2521]) begin
            regVec_2521 <= _zz_regVec_0;
          end
          if(_zz_1[2522]) begin
            regVec_2522 <= _zz_regVec_0;
          end
          if(_zz_1[2523]) begin
            regVec_2523 <= _zz_regVec_0;
          end
          if(_zz_1[2524]) begin
            regVec_2524 <= _zz_regVec_0;
          end
          if(_zz_1[2525]) begin
            regVec_2525 <= _zz_regVec_0;
          end
          if(_zz_1[2526]) begin
            regVec_2526 <= _zz_regVec_0;
          end
          if(_zz_1[2527]) begin
            regVec_2527 <= _zz_regVec_0;
          end
          if(_zz_1[2528]) begin
            regVec_2528 <= _zz_regVec_0;
          end
          if(_zz_1[2529]) begin
            regVec_2529 <= _zz_regVec_0;
          end
          if(_zz_1[2530]) begin
            regVec_2530 <= _zz_regVec_0;
          end
          if(_zz_1[2531]) begin
            regVec_2531 <= _zz_regVec_0;
          end
          if(_zz_1[2532]) begin
            regVec_2532 <= _zz_regVec_0;
          end
          if(_zz_1[2533]) begin
            regVec_2533 <= _zz_regVec_0;
          end
          if(_zz_1[2534]) begin
            regVec_2534 <= _zz_regVec_0;
          end
          if(_zz_1[2535]) begin
            regVec_2535 <= _zz_regVec_0;
          end
          if(_zz_1[2536]) begin
            regVec_2536 <= _zz_regVec_0;
          end
          if(_zz_1[2537]) begin
            regVec_2537 <= _zz_regVec_0;
          end
          if(_zz_1[2538]) begin
            regVec_2538 <= _zz_regVec_0;
          end
          if(_zz_1[2539]) begin
            regVec_2539 <= _zz_regVec_0;
          end
          if(_zz_1[2540]) begin
            regVec_2540 <= _zz_regVec_0;
          end
          if(_zz_1[2541]) begin
            regVec_2541 <= _zz_regVec_0;
          end
          if(_zz_1[2542]) begin
            regVec_2542 <= _zz_regVec_0;
          end
          if(_zz_1[2543]) begin
            regVec_2543 <= _zz_regVec_0;
          end
          if(_zz_1[2544]) begin
            regVec_2544 <= _zz_regVec_0;
          end
          if(_zz_1[2545]) begin
            regVec_2545 <= _zz_regVec_0;
          end
          if(_zz_1[2546]) begin
            regVec_2546 <= _zz_regVec_0;
          end
          if(_zz_1[2547]) begin
            regVec_2547 <= _zz_regVec_0;
          end
          if(_zz_1[2548]) begin
            regVec_2548 <= _zz_regVec_0;
          end
          if(_zz_1[2549]) begin
            regVec_2549 <= _zz_regVec_0;
          end
          if(_zz_1[2550]) begin
            regVec_2550 <= _zz_regVec_0;
          end
          if(_zz_1[2551]) begin
            regVec_2551 <= _zz_regVec_0;
          end
          if(_zz_1[2552]) begin
            regVec_2552 <= _zz_regVec_0;
          end
          if(_zz_1[2553]) begin
            regVec_2553 <= _zz_regVec_0;
          end
          if(_zz_1[2554]) begin
            regVec_2554 <= _zz_regVec_0;
          end
          if(_zz_1[2555]) begin
            regVec_2555 <= _zz_regVec_0;
          end
          if(_zz_1[2556]) begin
            regVec_2556 <= _zz_regVec_0;
          end
          if(_zz_1[2557]) begin
            regVec_2557 <= _zz_regVec_0;
          end
          if(_zz_1[2558]) begin
            regVec_2558 <= _zz_regVec_0;
          end
          if(_zz_1[2559]) begin
            regVec_2559 <= _zz_regVec_0;
          end
          if(_zz_1[2560]) begin
            regVec_2560 <= _zz_regVec_0;
          end
          if(_zz_1[2561]) begin
            regVec_2561 <= _zz_regVec_0;
          end
          if(_zz_1[2562]) begin
            regVec_2562 <= _zz_regVec_0;
          end
          if(_zz_1[2563]) begin
            regVec_2563 <= _zz_regVec_0;
          end
          if(_zz_1[2564]) begin
            regVec_2564 <= _zz_regVec_0;
          end
          if(_zz_1[2565]) begin
            regVec_2565 <= _zz_regVec_0;
          end
          if(_zz_1[2566]) begin
            regVec_2566 <= _zz_regVec_0;
          end
          if(_zz_1[2567]) begin
            regVec_2567 <= _zz_regVec_0;
          end
          if(_zz_1[2568]) begin
            regVec_2568 <= _zz_regVec_0;
          end
          if(_zz_1[2569]) begin
            regVec_2569 <= _zz_regVec_0;
          end
          if(_zz_1[2570]) begin
            regVec_2570 <= _zz_regVec_0;
          end
          if(_zz_1[2571]) begin
            regVec_2571 <= _zz_regVec_0;
          end
          if(_zz_1[2572]) begin
            regVec_2572 <= _zz_regVec_0;
          end
          if(_zz_1[2573]) begin
            regVec_2573 <= _zz_regVec_0;
          end
          if(_zz_1[2574]) begin
            regVec_2574 <= _zz_regVec_0;
          end
          if(_zz_1[2575]) begin
            regVec_2575 <= _zz_regVec_0;
          end
          if(_zz_1[2576]) begin
            regVec_2576 <= _zz_regVec_0;
          end
          if(_zz_1[2577]) begin
            regVec_2577 <= _zz_regVec_0;
          end
          if(_zz_1[2578]) begin
            regVec_2578 <= _zz_regVec_0;
          end
          if(_zz_1[2579]) begin
            regVec_2579 <= _zz_regVec_0;
          end
          if(_zz_1[2580]) begin
            regVec_2580 <= _zz_regVec_0;
          end
          if(_zz_1[2581]) begin
            regVec_2581 <= _zz_regVec_0;
          end
          if(_zz_1[2582]) begin
            regVec_2582 <= _zz_regVec_0;
          end
          if(_zz_1[2583]) begin
            regVec_2583 <= _zz_regVec_0;
          end
          if(_zz_1[2584]) begin
            regVec_2584 <= _zz_regVec_0;
          end
          if(_zz_1[2585]) begin
            regVec_2585 <= _zz_regVec_0;
          end
          if(_zz_1[2586]) begin
            regVec_2586 <= _zz_regVec_0;
          end
          if(_zz_1[2587]) begin
            regVec_2587 <= _zz_regVec_0;
          end
          if(_zz_1[2588]) begin
            regVec_2588 <= _zz_regVec_0;
          end
          if(_zz_1[2589]) begin
            regVec_2589 <= _zz_regVec_0;
          end
          if(_zz_1[2590]) begin
            regVec_2590 <= _zz_regVec_0;
          end
          if(_zz_1[2591]) begin
            regVec_2591 <= _zz_regVec_0;
          end
          if(_zz_1[2592]) begin
            regVec_2592 <= _zz_regVec_0;
          end
          if(_zz_1[2593]) begin
            regVec_2593 <= _zz_regVec_0;
          end
          if(_zz_1[2594]) begin
            regVec_2594 <= _zz_regVec_0;
          end
          if(_zz_1[2595]) begin
            regVec_2595 <= _zz_regVec_0;
          end
          if(_zz_1[2596]) begin
            regVec_2596 <= _zz_regVec_0;
          end
          if(_zz_1[2597]) begin
            regVec_2597 <= _zz_regVec_0;
          end
          if(_zz_1[2598]) begin
            regVec_2598 <= _zz_regVec_0;
          end
          if(_zz_1[2599]) begin
            regVec_2599 <= _zz_regVec_0;
          end
          if(_zz_1[2600]) begin
            regVec_2600 <= _zz_regVec_0;
          end
          if(_zz_1[2601]) begin
            regVec_2601 <= _zz_regVec_0;
          end
          if(_zz_1[2602]) begin
            regVec_2602 <= _zz_regVec_0;
          end
          if(_zz_1[2603]) begin
            regVec_2603 <= _zz_regVec_0;
          end
          if(_zz_1[2604]) begin
            regVec_2604 <= _zz_regVec_0;
          end
          if(_zz_1[2605]) begin
            regVec_2605 <= _zz_regVec_0;
          end
          if(_zz_1[2606]) begin
            regVec_2606 <= _zz_regVec_0;
          end
          if(_zz_1[2607]) begin
            regVec_2607 <= _zz_regVec_0;
          end
          if(_zz_1[2608]) begin
            regVec_2608 <= _zz_regVec_0;
          end
          if(_zz_1[2609]) begin
            regVec_2609 <= _zz_regVec_0;
          end
          if(_zz_1[2610]) begin
            regVec_2610 <= _zz_regVec_0;
          end
          if(_zz_1[2611]) begin
            regVec_2611 <= _zz_regVec_0;
          end
          if(_zz_1[2612]) begin
            regVec_2612 <= _zz_regVec_0;
          end
          if(_zz_1[2613]) begin
            regVec_2613 <= _zz_regVec_0;
          end
          if(_zz_1[2614]) begin
            regVec_2614 <= _zz_regVec_0;
          end
          if(_zz_1[2615]) begin
            regVec_2615 <= _zz_regVec_0;
          end
          if(_zz_1[2616]) begin
            regVec_2616 <= _zz_regVec_0;
          end
          if(_zz_1[2617]) begin
            regVec_2617 <= _zz_regVec_0;
          end
          if(_zz_1[2618]) begin
            regVec_2618 <= _zz_regVec_0;
          end
          if(_zz_1[2619]) begin
            regVec_2619 <= _zz_regVec_0;
          end
          if(_zz_1[2620]) begin
            regVec_2620 <= _zz_regVec_0;
          end
          if(_zz_1[2621]) begin
            regVec_2621 <= _zz_regVec_0;
          end
          if(_zz_1[2622]) begin
            regVec_2622 <= _zz_regVec_0;
          end
          if(_zz_1[2623]) begin
            regVec_2623 <= _zz_regVec_0;
          end
          if(_zz_1[2624]) begin
            regVec_2624 <= _zz_regVec_0;
          end
          if(_zz_1[2625]) begin
            regVec_2625 <= _zz_regVec_0;
          end
          if(_zz_1[2626]) begin
            regVec_2626 <= _zz_regVec_0;
          end
          if(_zz_1[2627]) begin
            regVec_2627 <= _zz_regVec_0;
          end
          if(_zz_1[2628]) begin
            regVec_2628 <= _zz_regVec_0;
          end
          if(_zz_1[2629]) begin
            regVec_2629 <= _zz_regVec_0;
          end
          if(_zz_1[2630]) begin
            regVec_2630 <= _zz_regVec_0;
          end
          if(_zz_1[2631]) begin
            regVec_2631 <= _zz_regVec_0;
          end
          if(_zz_1[2632]) begin
            regVec_2632 <= _zz_regVec_0;
          end
          if(_zz_1[2633]) begin
            regVec_2633 <= _zz_regVec_0;
          end
          if(_zz_1[2634]) begin
            regVec_2634 <= _zz_regVec_0;
          end
          if(_zz_1[2635]) begin
            regVec_2635 <= _zz_regVec_0;
          end
          if(_zz_1[2636]) begin
            regVec_2636 <= _zz_regVec_0;
          end
          if(_zz_1[2637]) begin
            regVec_2637 <= _zz_regVec_0;
          end
          if(_zz_1[2638]) begin
            regVec_2638 <= _zz_regVec_0;
          end
          if(_zz_1[2639]) begin
            regVec_2639 <= _zz_regVec_0;
          end
          if(_zz_1[2640]) begin
            regVec_2640 <= _zz_regVec_0;
          end
          if(_zz_1[2641]) begin
            regVec_2641 <= _zz_regVec_0;
          end
          if(_zz_1[2642]) begin
            regVec_2642 <= _zz_regVec_0;
          end
          if(_zz_1[2643]) begin
            regVec_2643 <= _zz_regVec_0;
          end
          if(_zz_1[2644]) begin
            regVec_2644 <= _zz_regVec_0;
          end
          if(_zz_1[2645]) begin
            regVec_2645 <= _zz_regVec_0;
          end
          if(_zz_1[2646]) begin
            regVec_2646 <= _zz_regVec_0;
          end
          if(_zz_1[2647]) begin
            regVec_2647 <= _zz_regVec_0;
          end
          if(_zz_1[2648]) begin
            regVec_2648 <= _zz_regVec_0;
          end
          if(_zz_1[2649]) begin
            regVec_2649 <= _zz_regVec_0;
          end
          if(_zz_1[2650]) begin
            regVec_2650 <= _zz_regVec_0;
          end
          if(_zz_1[2651]) begin
            regVec_2651 <= _zz_regVec_0;
          end
          if(_zz_1[2652]) begin
            regVec_2652 <= _zz_regVec_0;
          end
          if(_zz_1[2653]) begin
            regVec_2653 <= _zz_regVec_0;
          end
          if(_zz_1[2654]) begin
            regVec_2654 <= _zz_regVec_0;
          end
          if(_zz_1[2655]) begin
            regVec_2655 <= _zz_regVec_0;
          end
          if(_zz_1[2656]) begin
            regVec_2656 <= _zz_regVec_0;
          end
          if(_zz_1[2657]) begin
            regVec_2657 <= _zz_regVec_0;
          end
          if(_zz_1[2658]) begin
            regVec_2658 <= _zz_regVec_0;
          end
          if(_zz_1[2659]) begin
            regVec_2659 <= _zz_regVec_0;
          end
          if(_zz_1[2660]) begin
            regVec_2660 <= _zz_regVec_0;
          end
          if(_zz_1[2661]) begin
            regVec_2661 <= _zz_regVec_0;
          end
          if(_zz_1[2662]) begin
            regVec_2662 <= _zz_regVec_0;
          end
          if(_zz_1[2663]) begin
            regVec_2663 <= _zz_regVec_0;
          end
          if(_zz_1[2664]) begin
            regVec_2664 <= _zz_regVec_0;
          end
          if(_zz_1[2665]) begin
            regVec_2665 <= _zz_regVec_0;
          end
          if(_zz_1[2666]) begin
            regVec_2666 <= _zz_regVec_0;
          end
          if(_zz_1[2667]) begin
            regVec_2667 <= _zz_regVec_0;
          end
          if(_zz_1[2668]) begin
            regVec_2668 <= _zz_regVec_0;
          end
          if(_zz_1[2669]) begin
            regVec_2669 <= _zz_regVec_0;
          end
          if(_zz_1[2670]) begin
            regVec_2670 <= _zz_regVec_0;
          end
          if(_zz_1[2671]) begin
            regVec_2671 <= _zz_regVec_0;
          end
          if(_zz_1[2672]) begin
            regVec_2672 <= _zz_regVec_0;
          end
          if(_zz_1[2673]) begin
            regVec_2673 <= _zz_regVec_0;
          end
          if(_zz_1[2674]) begin
            regVec_2674 <= _zz_regVec_0;
          end
          if(_zz_1[2675]) begin
            regVec_2675 <= _zz_regVec_0;
          end
          if(_zz_1[2676]) begin
            regVec_2676 <= _zz_regVec_0;
          end
          if(_zz_1[2677]) begin
            regVec_2677 <= _zz_regVec_0;
          end
          if(_zz_1[2678]) begin
            regVec_2678 <= _zz_regVec_0;
          end
          if(_zz_1[2679]) begin
            regVec_2679 <= _zz_regVec_0;
          end
          if(_zz_1[2680]) begin
            regVec_2680 <= _zz_regVec_0;
          end
          if(_zz_1[2681]) begin
            regVec_2681 <= _zz_regVec_0;
          end
          if(_zz_1[2682]) begin
            regVec_2682 <= _zz_regVec_0;
          end
          if(_zz_1[2683]) begin
            regVec_2683 <= _zz_regVec_0;
          end
          if(_zz_1[2684]) begin
            regVec_2684 <= _zz_regVec_0;
          end
          if(_zz_1[2685]) begin
            regVec_2685 <= _zz_regVec_0;
          end
          if(_zz_1[2686]) begin
            regVec_2686 <= _zz_regVec_0;
          end
          if(_zz_1[2687]) begin
            regVec_2687 <= _zz_regVec_0;
          end
          if(_zz_1[2688]) begin
            regVec_2688 <= _zz_regVec_0;
          end
          if(_zz_1[2689]) begin
            regVec_2689 <= _zz_regVec_0;
          end
          if(_zz_1[2690]) begin
            regVec_2690 <= _zz_regVec_0;
          end
          if(_zz_1[2691]) begin
            regVec_2691 <= _zz_regVec_0;
          end
          if(_zz_1[2692]) begin
            regVec_2692 <= _zz_regVec_0;
          end
          if(_zz_1[2693]) begin
            regVec_2693 <= _zz_regVec_0;
          end
          if(_zz_1[2694]) begin
            regVec_2694 <= _zz_regVec_0;
          end
          if(_zz_1[2695]) begin
            regVec_2695 <= _zz_regVec_0;
          end
          if(_zz_1[2696]) begin
            regVec_2696 <= _zz_regVec_0;
          end
          if(_zz_1[2697]) begin
            regVec_2697 <= _zz_regVec_0;
          end
          if(_zz_1[2698]) begin
            regVec_2698 <= _zz_regVec_0;
          end
          if(_zz_1[2699]) begin
            regVec_2699 <= _zz_regVec_0;
          end
          if(_zz_1[2700]) begin
            regVec_2700 <= _zz_regVec_0;
          end
          if(_zz_1[2701]) begin
            regVec_2701 <= _zz_regVec_0;
          end
          if(_zz_1[2702]) begin
            regVec_2702 <= _zz_regVec_0;
          end
          if(_zz_1[2703]) begin
            regVec_2703 <= _zz_regVec_0;
          end
          if(_zz_1[2704]) begin
            regVec_2704 <= _zz_regVec_0;
          end
          if(_zz_1[2705]) begin
            regVec_2705 <= _zz_regVec_0;
          end
          if(_zz_1[2706]) begin
            regVec_2706 <= _zz_regVec_0;
          end
          if(_zz_1[2707]) begin
            regVec_2707 <= _zz_regVec_0;
          end
          if(_zz_1[2708]) begin
            regVec_2708 <= _zz_regVec_0;
          end
          if(_zz_1[2709]) begin
            regVec_2709 <= _zz_regVec_0;
          end
          if(_zz_1[2710]) begin
            regVec_2710 <= _zz_regVec_0;
          end
          if(_zz_1[2711]) begin
            regVec_2711 <= _zz_regVec_0;
          end
          if(_zz_1[2712]) begin
            regVec_2712 <= _zz_regVec_0;
          end
          if(_zz_1[2713]) begin
            regVec_2713 <= _zz_regVec_0;
          end
          if(_zz_1[2714]) begin
            regVec_2714 <= _zz_regVec_0;
          end
          if(_zz_1[2715]) begin
            regVec_2715 <= _zz_regVec_0;
          end
          if(_zz_1[2716]) begin
            regVec_2716 <= _zz_regVec_0;
          end
          if(_zz_1[2717]) begin
            regVec_2717 <= _zz_regVec_0;
          end
          if(_zz_1[2718]) begin
            regVec_2718 <= _zz_regVec_0;
          end
          if(_zz_1[2719]) begin
            regVec_2719 <= _zz_regVec_0;
          end
          if(_zz_1[2720]) begin
            regVec_2720 <= _zz_regVec_0;
          end
          if(_zz_1[2721]) begin
            regVec_2721 <= _zz_regVec_0;
          end
          if(_zz_1[2722]) begin
            regVec_2722 <= _zz_regVec_0;
          end
          if(_zz_1[2723]) begin
            regVec_2723 <= _zz_regVec_0;
          end
          if(_zz_1[2724]) begin
            regVec_2724 <= _zz_regVec_0;
          end
          if(_zz_1[2725]) begin
            regVec_2725 <= _zz_regVec_0;
          end
          if(_zz_1[2726]) begin
            regVec_2726 <= _zz_regVec_0;
          end
          if(_zz_1[2727]) begin
            regVec_2727 <= _zz_regVec_0;
          end
          if(_zz_1[2728]) begin
            regVec_2728 <= _zz_regVec_0;
          end
          if(_zz_1[2729]) begin
            regVec_2729 <= _zz_regVec_0;
          end
          if(_zz_1[2730]) begin
            regVec_2730 <= _zz_regVec_0;
          end
          if(_zz_1[2731]) begin
            regVec_2731 <= _zz_regVec_0;
          end
          if(_zz_1[2732]) begin
            regVec_2732 <= _zz_regVec_0;
          end
          if(_zz_1[2733]) begin
            regVec_2733 <= _zz_regVec_0;
          end
          if(_zz_1[2734]) begin
            regVec_2734 <= _zz_regVec_0;
          end
          if(_zz_1[2735]) begin
            regVec_2735 <= _zz_regVec_0;
          end
          if(_zz_1[2736]) begin
            regVec_2736 <= _zz_regVec_0;
          end
          if(_zz_1[2737]) begin
            regVec_2737 <= _zz_regVec_0;
          end
          if(_zz_1[2738]) begin
            regVec_2738 <= _zz_regVec_0;
          end
          if(_zz_1[2739]) begin
            regVec_2739 <= _zz_regVec_0;
          end
          if(_zz_1[2740]) begin
            regVec_2740 <= _zz_regVec_0;
          end
          if(_zz_1[2741]) begin
            regVec_2741 <= _zz_regVec_0;
          end
          if(_zz_1[2742]) begin
            regVec_2742 <= _zz_regVec_0;
          end
          if(_zz_1[2743]) begin
            regVec_2743 <= _zz_regVec_0;
          end
          if(_zz_1[2744]) begin
            regVec_2744 <= _zz_regVec_0;
          end
          if(_zz_1[2745]) begin
            regVec_2745 <= _zz_regVec_0;
          end
          if(_zz_1[2746]) begin
            regVec_2746 <= _zz_regVec_0;
          end
          if(_zz_1[2747]) begin
            regVec_2747 <= _zz_regVec_0;
          end
          if(_zz_1[2748]) begin
            regVec_2748 <= _zz_regVec_0;
          end
          if(_zz_1[2749]) begin
            regVec_2749 <= _zz_regVec_0;
          end
          if(_zz_1[2750]) begin
            regVec_2750 <= _zz_regVec_0;
          end
          if(_zz_1[2751]) begin
            regVec_2751 <= _zz_regVec_0;
          end
          if(_zz_1[2752]) begin
            regVec_2752 <= _zz_regVec_0;
          end
          if(_zz_1[2753]) begin
            regVec_2753 <= _zz_regVec_0;
          end
          if(_zz_1[2754]) begin
            regVec_2754 <= _zz_regVec_0;
          end
          if(_zz_1[2755]) begin
            regVec_2755 <= _zz_regVec_0;
          end
          if(_zz_1[2756]) begin
            regVec_2756 <= _zz_regVec_0;
          end
          if(_zz_1[2757]) begin
            regVec_2757 <= _zz_regVec_0;
          end
          if(_zz_1[2758]) begin
            regVec_2758 <= _zz_regVec_0;
          end
          if(_zz_1[2759]) begin
            regVec_2759 <= _zz_regVec_0;
          end
          if(_zz_1[2760]) begin
            regVec_2760 <= _zz_regVec_0;
          end
          if(_zz_1[2761]) begin
            regVec_2761 <= _zz_regVec_0;
          end
          if(_zz_1[2762]) begin
            regVec_2762 <= _zz_regVec_0;
          end
          if(_zz_1[2763]) begin
            regVec_2763 <= _zz_regVec_0;
          end
          if(_zz_1[2764]) begin
            regVec_2764 <= _zz_regVec_0;
          end
          if(_zz_1[2765]) begin
            regVec_2765 <= _zz_regVec_0;
          end
          if(_zz_1[2766]) begin
            regVec_2766 <= _zz_regVec_0;
          end
          if(_zz_1[2767]) begin
            regVec_2767 <= _zz_regVec_0;
          end
          if(_zz_1[2768]) begin
            regVec_2768 <= _zz_regVec_0;
          end
          if(_zz_1[2769]) begin
            regVec_2769 <= _zz_regVec_0;
          end
          if(_zz_1[2770]) begin
            regVec_2770 <= _zz_regVec_0;
          end
          if(_zz_1[2771]) begin
            regVec_2771 <= _zz_regVec_0;
          end
          if(_zz_1[2772]) begin
            regVec_2772 <= _zz_regVec_0;
          end
          if(_zz_1[2773]) begin
            regVec_2773 <= _zz_regVec_0;
          end
          if(_zz_1[2774]) begin
            regVec_2774 <= _zz_regVec_0;
          end
          if(_zz_1[2775]) begin
            regVec_2775 <= _zz_regVec_0;
          end
          if(_zz_1[2776]) begin
            regVec_2776 <= _zz_regVec_0;
          end
          if(_zz_1[2777]) begin
            regVec_2777 <= _zz_regVec_0;
          end
          if(_zz_1[2778]) begin
            regVec_2778 <= _zz_regVec_0;
          end
          if(_zz_1[2779]) begin
            regVec_2779 <= _zz_regVec_0;
          end
          if(_zz_1[2780]) begin
            regVec_2780 <= _zz_regVec_0;
          end
          if(_zz_1[2781]) begin
            regVec_2781 <= _zz_regVec_0;
          end
          if(_zz_1[2782]) begin
            regVec_2782 <= _zz_regVec_0;
          end
          if(_zz_1[2783]) begin
            regVec_2783 <= _zz_regVec_0;
          end
          if(_zz_1[2784]) begin
            regVec_2784 <= _zz_regVec_0;
          end
          if(_zz_1[2785]) begin
            regVec_2785 <= _zz_regVec_0;
          end
          if(_zz_1[2786]) begin
            regVec_2786 <= _zz_regVec_0;
          end
          if(_zz_1[2787]) begin
            regVec_2787 <= _zz_regVec_0;
          end
          if(_zz_1[2788]) begin
            regVec_2788 <= _zz_regVec_0;
          end
          if(_zz_1[2789]) begin
            regVec_2789 <= _zz_regVec_0;
          end
          if(_zz_1[2790]) begin
            regVec_2790 <= _zz_regVec_0;
          end
          if(_zz_1[2791]) begin
            regVec_2791 <= _zz_regVec_0;
          end
          if(_zz_1[2792]) begin
            regVec_2792 <= _zz_regVec_0;
          end
          if(_zz_1[2793]) begin
            regVec_2793 <= _zz_regVec_0;
          end
          if(_zz_1[2794]) begin
            regVec_2794 <= _zz_regVec_0;
          end
          if(_zz_1[2795]) begin
            regVec_2795 <= _zz_regVec_0;
          end
          if(_zz_1[2796]) begin
            regVec_2796 <= _zz_regVec_0;
          end
          if(_zz_1[2797]) begin
            regVec_2797 <= _zz_regVec_0;
          end
          if(_zz_1[2798]) begin
            regVec_2798 <= _zz_regVec_0;
          end
          if(_zz_1[2799]) begin
            regVec_2799 <= _zz_regVec_0;
          end
          if(_zz_1[2800]) begin
            regVec_2800 <= _zz_regVec_0;
          end
          if(_zz_1[2801]) begin
            regVec_2801 <= _zz_regVec_0;
          end
          if(_zz_1[2802]) begin
            regVec_2802 <= _zz_regVec_0;
          end
          if(_zz_1[2803]) begin
            regVec_2803 <= _zz_regVec_0;
          end
          if(_zz_1[2804]) begin
            regVec_2804 <= _zz_regVec_0;
          end
          if(_zz_1[2805]) begin
            regVec_2805 <= _zz_regVec_0;
          end
          if(_zz_1[2806]) begin
            regVec_2806 <= _zz_regVec_0;
          end
          if(_zz_1[2807]) begin
            regVec_2807 <= _zz_regVec_0;
          end
          if(_zz_1[2808]) begin
            regVec_2808 <= _zz_regVec_0;
          end
          if(_zz_1[2809]) begin
            regVec_2809 <= _zz_regVec_0;
          end
          if(_zz_1[2810]) begin
            regVec_2810 <= _zz_regVec_0;
          end
          if(_zz_1[2811]) begin
            regVec_2811 <= _zz_regVec_0;
          end
          if(_zz_1[2812]) begin
            regVec_2812 <= _zz_regVec_0;
          end
          if(_zz_1[2813]) begin
            regVec_2813 <= _zz_regVec_0;
          end
          if(_zz_1[2814]) begin
            regVec_2814 <= _zz_regVec_0;
          end
          if(_zz_1[2815]) begin
            regVec_2815 <= _zz_regVec_0;
          end
          if(_zz_1[2816]) begin
            regVec_2816 <= _zz_regVec_0;
          end
          if(_zz_1[2817]) begin
            regVec_2817 <= _zz_regVec_0;
          end
          if(_zz_1[2818]) begin
            regVec_2818 <= _zz_regVec_0;
          end
          if(_zz_1[2819]) begin
            regVec_2819 <= _zz_regVec_0;
          end
          if(_zz_1[2820]) begin
            regVec_2820 <= _zz_regVec_0;
          end
          if(_zz_1[2821]) begin
            regVec_2821 <= _zz_regVec_0;
          end
          if(_zz_1[2822]) begin
            regVec_2822 <= _zz_regVec_0;
          end
          if(_zz_1[2823]) begin
            regVec_2823 <= _zz_regVec_0;
          end
          if(_zz_1[2824]) begin
            regVec_2824 <= _zz_regVec_0;
          end
          if(_zz_1[2825]) begin
            regVec_2825 <= _zz_regVec_0;
          end
          if(_zz_1[2826]) begin
            regVec_2826 <= _zz_regVec_0;
          end
          if(_zz_1[2827]) begin
            regVec_2827 <= _zz_regVec_0;
          end
          if(_zz_1[2828]) begin
            regVec_2828 <= _zz_regVec_0;
          end
          if(_zz_1[2829]) begin
            regVec_2829 <= _zz_regVec_0;
          end
          if(_zz_1[2830]) begin
            regVec_2830 <= _zz_regVec_0;
          end
          if(_zz_1[2831]) begin
            regVec_2831 <= _zz_regVec_0;
          end
          if(_zz_1[2832]) begin
            regVec_2832 <= _zz_regVec_0;
          end
          if(_zz_1[2833]) begin
            regVec_2833 <= _zz_regVec_0;
          end
          if(_zz_1[2834]) begin
            regVec_2834 <= _zz_regVec_0;
          end
          if(_zz_1[2835]) begin
            regVec_2835 <= _zz_regVec_0;
          end
          if(_zz_1[2836]) begin
            regVec_2836 <= _zz_regVec_0;
          end
          if(_zz_1[2837]) begin
            regVec_2837 <= _zz_regVec_0;
          end
          if(_zz_1[2838]) begin
            regVec_2838 <= _zz_regVec_0;
          end
          if(_zz_1[2839]) begin
            regVec_2839 <= _zz_regVec_0;
          end
          if(_zz_1[2840]) begin
            regVec_2840 <= _zz_regVec_0;
          end
          if(_zz_1[2841]) begin
            regVec_2841 <= _zz_regVec_0;
          end
          if(_zz_1[2842]) begin
            regVec_2842 <= _zz_regVec_0;
          end
          if(_zz_1[2843]) begin
            regVec_2843 <= _zz_regVec_0;
          end
          if(_zz_1[2844]) begin
            regVec_2844 <= _zz_regVec_0;
          end
          if(_zz_1[2845]) begin
            regVec_2845 <= _zz_regVec_0;
          end
          if(_zz_1[2846]) begin
            regVec_2846 <= _zz_regVec_0;
          end
          if(_zz_1[2847]) begin
            regVec_2847 <= _zz_regVec_0;
          end
          if(_zz_1[2848]) begin
            regVec_2848 <= _zz_regVec_0;
          end
          if(_zz_1[2849]) begin
            regVec_2849 <= _zz_regVec_0;
          end
          if(_zz_1[2850]) begin
            regVec_2850 <= _zz_regVec_0;
          end
          if(_zz_1[2851]) begin
            regVec_2851 <= _zz_regVec_0;
          end
          if(_zz_1[2852]) begin
            regVec_2852 <= _zz_regVec_0;
          end
          if(_zz_1[2853]) begin
            regVec_2853 <= _zz_regVec_0;
          end
          if(_zz_1[2854]) begin
            regVec_2854 <= _zz_regVec_0;
          end
          if(_zz_1[2855]) begin
            regVec_2855 <= _zz_regVec_0;
          end
          if(_zz_1[2856]) begin
            regVec_2856 <= _zz_regVec_0;
          end
          if(_zz_1[2857]) begin
            regVec_2857 <= _zz_regVec_0;
          end
          if(_zz_1[2858]) begin
            regVec_2858 <= _zz_regVec_0;
          end
          if(_zz_1[2859]) begin
            regVec_2859 <= _zz_regVec_0;
          end
          if(_zz_1[2860]) begin
            regVec_2860 <= _zz_regVec_0;
          end
          if(_zz_1[2861]) begin
            regVec_2861 <= _zz_regVec_0;
          end
          if(_zz_1[2862]) begin
            regVec_2862 <= _zz_regVec_0;
          end
          if(_zz_1[2863]) begin
            regVec_2863 <= _zz_regVec_0;
          end
          if(_zz_1[2864]) begin
            regVec_2864 <= _zz_regVec_0;
          end
          if(_zz_1[2865]) begin
            regVec_2865 <= _zz_regVec_0;
          end
          if(_zz_1[2866]) begin
            regVec_2866 <= _zz_regVec_0;
          end
          if(_zz_1[2867]) begin
            regVec_2867 <= _zz_regVec_0;
          end
          if(_zz_1[2868]) begin
            regVec_2868 <= _zz_regVec_0;
          end
          if(_zz_1[2869]) begin
            regVec_2869 <= _zz_regVec_0;
          end
          if(_zz_1[2870]) begin
            regVec_2870 <= _zz_regVec_0;
          end
          if(_zz_1[2871]) begin
            regVec_2871 <= _zz_regVec_0;
          end
          if(_zz_1[2872]) begin
            regVec_2872 <= _zz_regVec_0;
          end
          if(_zz_1[2873]) begin
            regVec_2873 <= _zz_regVec_0;
          end
          if(_zz_1[2874]) begin
            regVec_2874 <= _zz_regVec_0;
          end
          if(_zz_1[2875]) begin
            regVec_2875 <= _zz_regVec_0;
          end
          if(_zz_1[2876]) begin
            regVec_2876 <= _zz_regVec_0;
          end
          if(_zz_1[2877]) begin
            regVec_2877 <= _zz_regVec_0;
          end
          if(_zz_1[2878]) begin
            regVec_2878 <= _zz_regVec_0;
          end
          if(_zz_1[2879]) begin
            regVec_2879 <= _zz_regVec_0;
          end
          if(_zz_1[2880]) begin
            regVec_2880 <= _zz_regVec_0;
          end
          if(_zz_1[2881]) begin
            regVec_2881 <= _zz_regVec_0;
          end
          if(_zz_1[2882]) begin
            regVec_2882 <= _zz_regVec_0;
          end
          if(_zz_1[2883]) begin
            regVec_2883 <= _zz_regVec_0;
          end
          if(_zz_1[2884]) begin
            regVec_2884 <= _zz_regVec_0;
          end
          if(_zz_1[2885]) begin
            regVec_2885 <= _zz_regVec_0;
          end
          if(_zz_1[2886]) begin
            regVec_2886 <= _zz_regVec_0;
          end
          if(_zz_1[2887]) begin
            regVec_2887 <= _zz_regVec_0;
          end
          if(_zz_1[2888]) begin
            regVec_2888 <= _zz_regVec_0;
          end
          if(_zz_1[2889]) begin
            regVec_2889 <= _zz_regVec_0;
          end
          if(_zz_1[2890]) begin
            regVec_2890 <= _zz_regVec_0;
          end
          if(_zz_1[2891]) begin
            regVec_2891 <= _zz_regVec_0;
          end
          if(_zz_1[2892]) begin
            regVec_2892 <= _zz_regVec_0;
          end
          if(_zz_1[2893]) begin
            regVec_2893 <= _zz_regVec_0;
          end
          if(_zz_1[2894]) begin
            regVec_2894 <= _zz_regVec_0;
          end
          if(_zz_1[2895]) begin
            regVec_2895 <= _zz_regVec_0;
          end
          if(_zz_1[2896]) begin
            regVec_2896 <= _zz_regVec_0;
          end
          if(_zz_1[2897]) begin
            regVec_2897 <= _zz_regVec_0;
          end
          if(_zz_1[2898]) begin
            regVec_2898 <= _zz_regVec_0;
          end
          if(_zz_1[2899]) begin
            regVec_2899 <= _zz_regVec_0;
          end
          if(_zz_1[2900]) begin
            regVec_2900 <= _zz_regVec_0;
          end
          if(_zz_1[2901]) begin
            regVec_2901 <= _zz_regVec_0;
          end
          if(_zz_1[2902]) begin
            regVec_2902 <= _zz_regVec_0;
          end
          if(_zz_1[2903]) begin
            regVec_2903 <= _zz_regVec_0;
          end
          if(_zz_1[2904]) begin
            regVec_2904 <= _zz_regVec_0;
          end
          if(_zz_1[2905]) begin
            regVec_2905 <= _zz_regVec_0;
          end
          if(_zz_1[2906]) begin
            regVec_2906 <= _zz_regVec_0;
          end
          if(_zz_1[2907]) begin
            regVec_2907 <= _zz_regVec_0;
          end
          if(_zz_1[2908]) begin
            regVec_2908 <= _zz_regVec_0;
          end
          if(_zz_1[2909]) begin
            regVec_2909 <= _zz_regVec_0;
          end
          if(_zz_1[2910]) begin
            regVec_2910 <= _zz_regVec_0;
          end
          if(_zz_1[2911]) begin
            regVec_2911 <= _zz_regVec_0;
          end
          if(_zz_1[2912]) begin
            regVec_2912 <= _zz_regVec_0;
          end
          if(_zz_1[2913]) begin
            regVec_2913 <= _zz_regVec_0;
          end
          if(_zz_1[2914]) begin
            regVec_2914 <= _zz_regVec_0;
          end
          if(_zz_1[2915]) begin
            regVec_2915 <= _zz_regVec_0;
          end
          if(_zz_1[2916]) begin
            regVec_2916 <= _zz_regVec_0;
          end
          if(_zz_1[2917]) begin
            regVec_2917 <= _zz_regVec_0;
          end
          if(_zz_1[2918]) begin
            regVec_2918 <= _zz_regVec_0;
          end
          if(_zz_1[2919]) begin
            regVec_2919 <= _zz_regVec_0;
          end
          if(_zz_1[2920]) begin
            regVec_2920 <= _zz_regVec_0;
          end
          if(_zz_1[2921]) begin
            regVec_2921 <= _zz_regVec_0;
          end
          if(_zz_1[2922]) begin
            regVec_2922 <= _zz_regVec_0;
          end
          if(_zz_1[2923]) begin
            regVec_2923 <= _zz_regVec_0;
          end
          if(_zz_1[2924]) begin
            regVec_2924 <= _zz_regVec_0;
          end
          if(_zz_1[2925]) begin
            regVec_2925 <= _zz_regVec_0;
          end
          if(_zz_1[2926]) begin
            regVec_2926 <= _zz_regVec_0;
          end
          if(_zz_1[2927]) begin
            regVec_2927 <= _zz_regVec_0;
          end
          if(_zz_1[2928]) begin
            regVec_2928 <= _zz_regVec_0;
          end
          if(_zz_1[2929]) begin
            regVec_2929 <= _zz_regVec_0;
          end
          if(_zz_1[2930]) begin
            regVec_2930 <= _zz_regVec_0;
          end
          if(_zz_1[2931]) begin
            regVec_2931 <= _zz_regVec_0;
          end
          if(_zz_1[2932]) begin
            regVec_2932 <= _zz_regVec_0;
          end
          if(_zz_1[2933]) begin
            regVec_2933 <= _zz_regVec_0;
          end
          if(_zz_1[2934]) begin
            regVec_2934 <= _zz_regVec_0;
          end
          if(_zz_1[2935]) begin
            regVec_2935 <= _zz_regVec_0;
          end
          if(_zz_1[2936]) begin
            regVec_2936 <= _zz_regVec_0;
          end
          if(_zz_1[2937]) begin
            regVec_2937 <= _zz_regVec_0;
          end
          if(_zz_1[2938]) begin
            regVec_2938 <= _zz_regVec_0;
          end
          if(_zz_1[2939]) begin
            regVec_2939 <= _zz_regVec_0;
          end
          if(_zz_1[2940]) begin
            regVec_2940 <= _zz_regVec_0;
          end
          if(_zz_1[2941]) begin
            regVec_2941 <= _zz_regVec_0;
          end
          if(_zz_1[2942]) begin
            regVec_2942 <= _zz_regVec_0;
          end
          if(_zz_1[2943]) begin
            regVec_2943 <= _zz_regVec_0;
          end
          if(_zz_1[2944]) begin
            regVec_2944 <= _zz_regVec_0;
          end
          if(_zz_1[2945]) begin
            regVec_2945 <= _zz_regVec_0;
          end
          if(_zz_1[2946]) begin
            regVec_2946 <= _zz_regVec_0;
          end
          if(_zz_1[2947]) begin
            regVec_2947 <= _zz_regVec_0;
          end
          if(_zz_1[2948]) begin
            regVec_2948 <= _zz_regVec_0;
          end
          if(_zz_1[2949]) begin
            regVec_2949 <= _zz_regVec_0;
          end
          if(_zz_1[2950]) begin
            regVec_2950 <= _zz_regVec_0;
          end
          if(_zz_1[2951]) begin
            regVec_2951 <= _zz_regVec_0;
          end
          if(_zz_1[2952]) begin
            regVec_2952 <= _zz_regVec_0;
          end
          if(_zz_1[2953]) begin
            regVec_2953 <= _zz_regVec_0;
          end
          if(_zz_1[2954]) begin
            regVec_2954 <= _zz_regVec_0;
          end
          if(_zz_1[2955]) begin
            regVec_2955 <= _zz_regVec_0;
          end
          if(_zz_1[2956]) begin
            regVec_2956 <= _zz_regVec_0;
          end
          if(_zz_1[2957]) begin
            regVec_2957 <= _zz_regVec_0;
          end
          if(_zz_1[2958]) begin
            regVec_2958 <= _zz_regVec_0;
          end
          if(_zz_1[2959]) begin
            regVec_2959 <= _zz_regVec_0;
          end
          if(_zz_1[2960]) begin
            regVec_2960 <= _zz_regVec_0;
          end
          if(_zz_1[2961]) begin
            regVec_2961 <= _zz_regVec_0;
          end
          if(_zz_1[2962]) begin
            regVec_2962 <= _zz_regVec_0;
          end
          if(_zz_1[2963]) begin
            regVec_2963 <= _zz_regVec_0;
          end
          if(_zz_1[2964]) begin
            regVec_2964 <= _zz_regVec_0;
          end
          if(_zz_1[2965]) begin
            regVec_2965 <= _zz_regVec_0;
          end
          if(_zz_1[2966]) begin
            regVec_2966 <= _zz_regVec_0;
          end
          if(_zz_1[2967]) begin
            regVec_2967 <= _zz_regVec_0;
          end
          if(_zz_1[2968]) begin
            regVec_2968 <= _zz_regVec_0;
          end
          if(_zz_1[2969]) begin
            regVec_2969 <= _zz_regVec_0;
          end
          if(_zz_1[2970]) begin
            regVec_2970 <= _zz_regVec_0;
          end
          if(_zz_1[2971]) begin
            regVec_2971 <= _zz_regVec_0;
          end
          if(_zz_1[2972]) begin
            regVec_2972 <= _zz_regVec_0;
          end
          if(_zz_1[2973]) begin
            regVec_2973 <= _zz_regVec_0;
          end
          if(_zz_1[2974]) begin
            regVec_2974 <= _zz_regVec_0;
          end
          if(_zz_1[2975]) begin
            regVec_2975 <= _zz_regVec_0;
          end
          if(_zz_1[2976]) begin
            regVec_2976 <= _zz_regVec_0;
          end
          if(_zz_1[2977]) begin
            regVec_2977 <= _zz_regVec_0;
          end
          if(_zz_1[2978]) begin
            regVec_2978 <= _zz_regVec_0;
          end
          if(_zz_1[2979]) begin
            regVec_2979 <= _zz_regVec_0;
          end
          if(_zz_1[2980]) begin
            regVec_2980 <= _zz_regVec_0;
          end
          if(_zz_1[2981]) begin
            regVec_2981 <= _zz_regVec_0;
          end
          if(_zz_1[2982]) begin
            regVec_2982 <= _zz_regVec_0;
          end
          if(_zz_1[2983]) begin
            regVec_2983 <= _zz_regVec_0;
          end
          if(_zz_1[2984]) begin
            regVec_2984 <= _zz_regVec_0;
          end
          if(_zz_1[2985]) begin
            regVec_2985 <= _zz_regVec_0;
          end
          if(_zz_1[2986]) begin
            regVec_2986 <= _zz_regVec_0;
          end
          if(_zz_1[2987]) begin
            regVec_2987 <= _zz_regVec_0;
          end
          if(_zz_1[2988]) begin
            regVec_2988 <= _zz_regVec_0;
          end
          if(_zz_1[2989]) begin
            regVec_2989 <= _zz_regVec_0;
          end
          if(_zz_1[2990]) begin
            regVec_2990 <= _zz_regVec_0;
          end
          if(_zz_1[2991]) begin
            regVec_2991 <= _zz_regVec_0;
          end
          if(_zz_1[2992]) begin
            regVec_2992 <= _zz_regVec_0;
          end
          if(_zz_1[2993]) begin
            regVec_2993 <= _zz_regVec_0;
          end
          if(_zz_1[2994]) begin
            regVec_2994 <= _zz_regVec_0;
          end
          if(_zz_1[2995]) begin
            regVec_2995 <= _zz_regVec_0;
          end
          if(_zz_1[2996]) begin
            regVec_2996 <= _zz_regVec_0;
          end
          if(_zz_1[2997]) begin
            regVec_2997 <= _zz_regVec_0;
          end
          if(_zz_1[2998]) begin
            regVec_2998 <= _zz_regVec_0;
          end
          if(_zz_1[2999]) begin
            regVec_2999 <= _zz_regVec_0;
          end
          if(_zz_1[3000]) begin
            regVec_3000 <= _zz_regVec_0;
          end
          if(_zz_1[3001]) begin
            regVec_3001 <= _zz_regVec_0;
          end
          if(_zz_1[3002]) begin
            regVec_3002 <= _zz_regVec_0;
          end
          if(_zz_1[3003]) begin
            regVec_3003 <= _zz_regVec_0;
          end
          if(_zz_1[3004]) begin
            regVec_3004 <= _zz_regVec_0;
          end
          if(_zz_1[3005]) begin
            regVec_3005 <= _zz_regVec_0;
          end
          if(_zz_1[3006]) begin
            regVec_3006 <= _zz_regVec_0;
          end
          if(_zz_1[3007]) begin
            regVec_3007 <= _zz_regVec_0;
          end
          if(_zz_1[3008]) begin
            regVec_3008 <= _zz_regVec_0;
          end
          if(_zz_1[3009]) begin
            regVec_3009 <= _zz_regVec_0;
          end
          if(_zz_1[3010]) begin
            regVec_3010 <= _zz_regVec_0;
          end
          if(_zz_1[3011]) begin
            regVec_3011 <= _zz_regVec_0;
          end
          if(_zz_1[3012]) begin
            regVec_3012 <= _zz_regVec_0;
          end
          if(_zz_1[3013]) begin
            regVec_3013 <= _zz_regVec_0;
          end
          if(_zz_1[3014]) begin
            regVec_3014 <= _zz_regVec_0;
          end
          if(_zz_1[3015]) begin
            regVec_3015 <= _zz_regVec_0;
          end
          if(_zz_1[3016]) begin
            regVec_3016 <= _zz_regVec_0;
          end
          if(_zz_1[3017]) begin
            regVec_3017 <= _zz_regVec_0;
          end
          if(_zz_1[3018]) begin
            regVec_3018 <= _zz_regVec_0;
          end
          if(_zz_1[3019]) begin
            regVec_3019 <= _zz_regVec_0;
          end
          if(_zz_1[3020]) begin
            regVec_3020 <= _zz_regVec_0;
          end
          if(_zz_1[3021]) begin
            regVec_3021 <= _zz_regVec_0;
          end
          if(_zz_1[3022]) begin
            regVec_3022 <= _zz_regVec_0;
          end
          if(_zz_1[3023]) begin
            regVec_3023 <= _zz_regVec_0;
          end
          if(_zz_1[3024]) begin
            regVec_3024 <= _zz_regVec_0;
          end
          if(_zz_1[3025]) begin
            regVec_3025 <= _zz_regVec_0;
          end
          if(_zz_1[3026]) begin
            regVec_3026 <= _zz_regVec_0;
          end
          if(_zz_1[3027]) begin
            regVec_3027 <= _zz_regVec_0;
          end
          if(_zz_1[3028]) begin
            regVec_3028 <= _zz_regVec_0;
          end
          if(_zz_1[3029]) begin
            regVec_3029 <= _zz_regVec_0;
          end
          if(_zz_1[3030]) begin
            regVec_3030 <= _zz_regVec_0;
          end
          if(_zz_1[3031]) begin
            regVec_3031 <= _zz_regVec_0;
          end
          if(_zz_1[3032]) begin
            regVec_3032 <= _zz_regVec_0;
          end
          if(_zz_1[3033]) begin
            regVec_3033 <= _zz_regVec_0;
          end
          if(_zz_1[3034]) begin
            regVec_3034 <= _zz_regVec_0;
          end
          if(_zz_1[3035]) begin
            regVec_3035 <= _zz_regVec_0;
          end
          if(_zz_1[3036]) begin
            regVec_3036 <= _zz_regVec_0;
          end
          if(_zz_1[3037]) begin
            regVec_3037 <= _zz_regVec_0;
          end
          if(_zz_1[3038]) begin
            regVec_3038 <= _zz_regVec_0;
          end
          if(_zz_1[3039]) begin
            regVec_3039 <= _zz_regVec_0;
          end
          if(_zz_1[3040]) begin
            regVec_3040 <= _zz_regVec_0;
          end
          if(_zz_1[3041]) begin
            regVec_3041 <= _zz_regVec_0;
          end
          if(_zz_1[3042]) begin
            regVec_3042 <= _zz_regVec_0;
          end
          if(_zz_1[3043]) begin
            regVec_3043 <= _zz_regVec_0;
          end
          if(_zz_1[3044]) begin
            regVec_3044 <= _zz_regVec_0;
          end
          if(_zz_1[3045]) begin
            regVec_3045 <= _zz_regVec_0;
          end
          if(_zz_1[3046]) begin
            regVec_3046 <= _zz_regVec_0;
          end
          if(_zz_1[3047]) begin
            regVec_3047 <= _zz_regVec_0;
          end
          if(_zz_1[3048]) begin
            regVec_3048 <= _zz_regVec_0;
          end
          if(_zz_1[3049]) begin
            regVec_3049 <= _zz_regVec_0;
          end
          if(_zz_1[3050]) begin
            regVec_3050 <= _zz_regVec_0;
          end
          if(_zz_1[3051]) begin
            regVec_3051 <= _zz_regVec_0;
          end
          if(_zz_1[3052]) begin
            regVec_3052 <= _zz_regVec_0;
          end
          if(_zz_1[3053]) begin
            regVec_3053 <= _zz_regVec_0;
          end
          if(_zz_1[3054]) begin
            regVec_3054 <= _zz_regVec_0;
          end
          if(_zz_1[3055]) begin
            regVec_3055 <= _zz_regVec_0;
          end
          if(_zz_1[3056]) begin
            regVec_3056 <= _zz_regVec_0;
          end
          if(_zz_1[3057]) begin
            regVec_3057 <= _zz_regVec_0;
          end
          if(_zz_1[3058]) begin
            regVec_3058 <= _zz_regVec_0;
          end
          if(_zz_1[3059]) begin
            regVec_3059 <= _zz_regVec_0;
          end
          if(_zz_1[3060]) begin
            regVec_3060 <= _zz_regVec_0;
          end
          if(_zz_1[3061]) begin
            regVec_3061 <= _zz_regVec_0;
          end
          if(_zz_1[3062]) begin
            regVec_3062 <= _zz_regVec_0;
          end
          if(_zz_1[3063]) begin
            regVec_3063 <= _zz_regVec_0;
          end
          if(_zz_1[3064]) begin
            regVec_3064 <= _zz_regVec_0;
          end
          if(_zz_1[3065]) begin
            regVec_3065 <= _zz_regVec_0;
          end
          if(_zz_1[3066]) begin
            regVec_3066 <= _zz_regVec_0;
          end
          if(_zz_1[3067]) begin
            regVec_3067 <= _zz_regVec_0;
          end
          if(_zz_1[3068]) begin
            regVec_3068 <= _zz_regVec_0;
          end
          if(_zz_1[3069]) begin
            regVec_3069 <= _zz_regVec_0;
          end
          if(_zz_1[3070]) begin
            regVec_3070 <= _zz_regVec_0;
          end
          if(_zz_1[3071]) begin
            regVec_3071 <= _zz_regVec_0;
          end
          if(_zz_1[3072]) begin
            regVec_3072 <= _zz_regVec_0;
          end
          if(_zz_1[3073]) begin
            regVec_3073 <= _zz_regVec_0;
          end
          if(_zz_1[3074]) begin
            regVec_3074 <= _zz_regVec_0;
          end
          if(_zz_1[3075]) begin
            regVec_3075 <= _zz_regVec_0;
          end
          if(_zz_1[3076]) begin
            regVec_3076 <= _zz_regVec_0;
          end
          if(_zz_1[3077]) begin
            regVec_3077 <= _zz_regVec_0;
          end
          if(_zz_1[3078]) begin
            regVec_3078 <= _zz_regVec_0;
          end
          if(_zz_1[3079]) begin
            regVec_3079 <= _zz_regVec_0;
          end
          if(_zz_1[3080]) begin
            regVec_3080 <= _zz_regVec_0;
          end
          if(_zz_1[3081]) begin
            regVec_3081 <= _zz_regVec_0;
          end
          if(_zz_1[3082]) begin
            regVec_3082 <= _zz_regVec_0;
          end
          if(_zz_1[3083]) begin
            regVec_3083 <= _zz_regVec_0;
          end
          if(_zz_1[3084]) begin
            regVec_3084 <= _zz_regVec_0;
          end
          if(_zz_1[3085]) begin
            regVec_3085 <= _zz_regVec_0;
          end
          if(_zz_1[3086]) begin
            regVec_3086 <= _zz_regVec_0;
          end
          if(_zz_1[3087]) begin
            regVec_3087 <= _zz_regVec_0;
          end
          if(_zz_1[3088]) begin
            regVec_3088 <= _zz_regVec_0;
          end
          if(_zz_1[3089]) begin
            regVec_3089 <= _zz_regVec_0;
          end
          if(_zz_1[3090]) begin
            regVec_3090 <= _zz_regVec_0;
          end
          if(_zz_1[3091]) begin
            regVec_3091 <= _zz_regVec_0;
          end
          if(_zz_1[3092]) begin
            regVec_3092 <= _zz_regVec_0;
          end
          if(_zz_1[3093]) begin
            regVec_3093 <= _zz_regVec_0;
          end
          if(_zz_1[3094]) begin
            regVec_3094 <= _zz_regVec_0;
          end
          if(_zz_1[3095]) begin
            regVec_3095 <= _zz_regVec_0;
          end
          if(_zz_1[3096]) begin
            regVec_3096 <= _zz_regVec_0;
          end
          if(_zz_1[3097]) begin
            regVec_3097 <= _zz_regVec_0;
          end
          if(_zz_1[3098]) begin
            regVec_3098 <= _zz_regVec_0;
          end
          if(_zz_1[3099]) begin
            regVec_3099 <= _zz_regVec_0;
          end
          if(_zz_1[3100]) begin
            regVec_3100 <= _zz_regVec_0;
          end
          if(_zz_1[3101]) begin
            regVec_3101 <= _zz_regVec_0;
          end
          if(_zz_1[3102]) begin
            regVec_3102 <= _zz_regVec_0;
          end
          if(_zz_1[3103]) begin
            regVec_3103 <= _zz_regVec_0;
          end
          if(_zz_1[3104]) begin
            regVec_3104 <= _zz_regVec_0;
          end
          if(_zz_1[3105]) begin
            regVec_3105 <= _zz_regVec_0;
          end
          if(_zz_1[3106]) begin
            regVec_3106 <= _zz_regVec_0;
          end
          if(_zz_1[3107]) begin
            regVec_3107 <= _zz_regVec_0;
          end
          if(_zz_1[3108]) begin
            regVec_3108 <= _zz_regVec_0;
          end
          if(_zz_1[3109]) begin
            regVec_3109 <= _zz_regVec_0;
          end
          if(_zz_1[3110]) begin
            regVec_3110 <= _zz_regVec_0;
          end
          if(_zz_1[3111]) begin
            regVec_3111 <= _zz_regVec_0;
          end
          if(_zz_1[3112]) begin
            regVec_3112 <= _zz_regVec_0;
          end
          if(_zz_1[3113]) begin
            regVec_3113 <= _zz_regVec_0;
          end
          if(_zz_1[3114]) begin
            regVec_3114 <= _zz_regVec_0;
          end
          if(_zz_1[3115]) begin
            regVec_3115 <= _zz_regVec_0;
          end
          if(_zz_1[3116]) begin
            regVec_3116 <= _zz_regVec_0;
          end
          if(_zz_1[3117]) begin
            regVec_3117 <= _zz_regVec_0;
          end
          if(_zz_1[3118]) begin
            regVec_3118 <= _zz_regVec_0;
          end
          if(_zz_1[3119]) begin
            regVec_3119 <= _zz_regVec_0;
          end
          if(_zz_1[3120]) begin
            regVec_3120 <= _zz_regVec_0;
          end
          if(_zz_1[3121]) begin
            regVec_3121 <= _zz_regVec_0;
          end
          if(_zz_1[3122]) begin
            regVec_3122 <= _zz_regVec_0;
          end
          if(_zz_1[3123]) begin
            regVec_3123 <= _zz_regVec_0;
          end
          if(_zz_1[3124]) begin
            regVec_3124 <= _zz_regVec_0;
          end
          if(_zz_1[3125]) begin
            regVec_3125 <= _zz_regVec_0;
          end
          if(_zz_1[3126]) begin
            regVec_3126 <= _zz_regVec_0;
          end
          if(_zz_1[3127]) begin
            regVec_3127 <= _zz_regVec_0;
          end
          if(_zz_1[3128]) begin
            regVec_3128 <= _zz_regVec_0;
          end
          if(_zz_1[3129]) begin
            regVec_3129 <= _zz_regVec_0;
          end
          if(_zz_1[3130]) begin
            regVec_3130 <= _zz_regVec_0;
          end
          if(_zz_1[3131]) begin
            regVec_3131 <= _zz_regVec_0;
          end
          if(_zz_1[3132]) begin
            regVec_3132 <= _zz_regVec_0;
          end
          if(_zz_1[3133]) begin
            regVec_3133 <= _zz_regVec_0;
          end
          if(_zz_1[3134]) begin
            regVec_3134 <= _zz_regVec_0;
          end
          if(_zz_1[3135]) begin
            regVec_3135 <= _zz_regVec_0;
          end
          if(_zz_1[3136]) begin
            regVec_3136 <= _zz_regVec_0;
          end
          if(_zz_1[3137]) begin
            regVec_3137 <= _zz_regVec_0;
          end
          if(_zz_1[3138]) begin
            regVec_3138 <= _zz_regVec_0;
          end
          if(_zz_1[3139]) begin
            regVec_3139 <= _zz_regVec_0;
          end
          if(_zz_1[3140]) begin
            regVec_3140 <= _zz_regVec_0;
          end
          if(_zz_1[3141]) begin
            regVec_3141 <= _zz_regVec_0;
          end
          if(_zz_1[3142]) begin
            regVec_3142 <= _zz_regVec_0;
          end
          if(_zz_1[3143]) begin
            regVec_3143 <= _zz_regVec_0;
          end
          if(_zz_1[3144]) begin
            regVec_3144 <= _zz_regVec_0;
          end
          if(_zz_1[3145]) begin
            regVec_3145 <= _zz_regVec_0;
          end
          if(_zz_1[3146]) begin
            regVec_3146 <= _zz_regVec_0;
          end
          if(_zz_1[3147]) begin
            regVec_3147 <= _zz_regVec_0;
          end
          if(_zz_1[3148]) begin
            regVec_3148 <= _zz_regVec_0;
          end
          if(_zz_1[3149]) begin
            regVec_3149 <= _zz_regVec_0;
          end
          if(_zz_1[3150]) begin
            regVec_3150 <= _zz_regVec_0;
          end
          if(_zz_1[3151]) begin
            regVec_3151 <= _zz_regVec_0;
          end
          if(_zz_1[3152]) begin
            regVec_3152 <= _zz_regVec_0;
          end
          if(_zz_1[3153]) begin
            regVec_3153 <= _zz_regVec_0;
          end
          if(_zz_1[3154]) begin
            regVec_3154 <= _zz_regVec_0;
          end
          if(_zz_1[3155]) begin
            regVec_3155 <= _zz_regVec_0;
          end
          if(_zz_1[3156]) begin
            regVec_3156 <= _zz_regVec_0;
          end
          if(_zz_1[3157]) begin
            regVec_3157 <= _zz_regVec_0;
          end
          if(_zz_1[3158]) begin
            regVec_3158 <= _zz_regVec_0;
          end
          if(_zz_1[3159]) begin
            regVec_3159 <= _zz_regVec_0;
          end
          if(_zz_1[3160]) begin
            regVec_3160 <= _zz_regVec_0;
          end
          if(_zz_1[3161]) begin
            regVec_3161 <= _zz_regVec_0;
          end
          if(_zz_1[3162]) begin
            regVec_3162 <= _zz_regVec_0;
          end
          if(_zz_1[3163]) begin
            regVec_3163 <= _zz_regVec_0;
          end
          if(_zz_1[3164]) begin
            regVec_3164 <= _zz_regVec_0;
          end
          if(_zz_1[3165]) begin
            regVec_3165 <= _zz_regVec_0;
          end
          if(_zz_1[3166]) begin
            regVec_3166 <= _zz_regVec_0;
          end
          if(_zz_1[3167]) begin
            regVec_3167 <= _zz_regVec_0;
          end
          if(_zz_1[3168]) begin
            regVec_3168 <= _zz_regVec_0;
          end
          if(_zz_1[3169]) begin
            regVec_3169 <= _zz_regVec_0;
          end
          if(_zz_1[3170]) begin
            regVec_3170 <= _zz_regVec_0;
          end
          if(_zz_1[3171]) begin
            regVec_3171 <= _zz_regVec_0;
          end
          if(_zz_1[3172]) begin
            regVec_3172 <= _zz_regVec_0;
          end
          if(_zz_1[3173]) begin
            regVec_3173 <= _zz_regVec_0;
          end
          if(_zz_1[3174]) begin
            regVec_3174 <= _zz_regVec_0;
          end
          if(_zz_1[3175]) begin
            regVec_3175 <= _zz_regVec_0;
          end
          if(_zz_1[3176]) begin
            regVec_3176 <= _zz_regVec_0;
          end
          if(_zz_1[3177]) begin
            regVec_3177 <= _zz_regVec_0;
          end
          if(_zz_1[3178]) begin
            regVec_3178 <= _zz_regVec_0;
          end
          if(_zz_1[3179]) begin
            regVec_3179 <= _zz_regVec_0;
          end
          if(_zz_1[3180]) begin
            regVec_3180 <= _zz_regVec_0;
          end
          if(_zz_1[3181]) begin
            regVec_3181 <= _zz_regVec_0;
          end
          if(_zz_1[3182]) begin
            regVec_3182 <= _zz_regVec_0;
          end
          if(_zz_1[3183]) begin
            regVec_3183 <= _zz_regVec_0;
          end
          if(_zz_1[3184]) begin
            regVec_3184 <= _zz_regVec_0;
          end
          if(_zz_1[3185]) begin
            regVec_3185 <= _zz_regVec_0;
          end
          if(_zz_1[3186]) begin
            regVec_3186 <= _zz_regVec_0;
          end
          if(_zz_1[3187]) begin
            regVec_3187 <= _zz_regVec_0;
          end
          if(_zz_1[3188]) begin
            regVec_3188 <= _zz_regVec_0;
          end
          if(_zz_1[3189]) begin
            regVec_3189 <= _zz_regVec_0;
          end
          if(_zz_1[3190]) begin
            regVec_3190 <= _zz_regVec_0;
          end
          if(_zz_1[3191]) begin
            regVec_3191 <= _zz_regVec_0;
          end
          if(_zz_1[3192]) begin
            regVec_3192 <= _zz_regVec_0;
          end
          if(_zz_1[3193]) begin
            regVec_3193 <= _zz_regVec_0;
          end
          if(_zz_1[3194]) begin
            regVec_3194 <= _zz_regVec_0;
          end
          if(_zz_1[3195]) begin
            regVec_3195 <= _zz_regVec_0;
          end
          if(_zz_1[3196]) begin
            regVec_3196 <= _zz_regVec_0;
          end
          if(_zz_1[3197]) begin
            regVec_3197 <= _zz_regVec_0;
          end
          if(_zz_1[3198]) begin
            regVec_3198 <= _zz_regVec_0;
          end
          if(_zz_1[3199]) begin
            regVec_3199 <= _zz_regVec_0;
          end
          if(_zz_1[3200]) begin
            regVec_3200 <= _zz_regVec_0;
          end
          if(_zz_1[3201]) begin
            regVec_3201 <= _zz_regVec_0;
          end
          if(_zz_1[3202]) begin
            regVec_3202 <= _zz_regVec_0;
          end
          if(_zz_1[3203]) begin
            regVec_3203 <= _zz_regVec_0;
          end
          if(_zz_1[3204]) begin
            regVec_3204 <= _zz_regVec_0;
          end
          if(_zz_1[3205]) begin
            regVec_3205 <= _zz_regVec_0;
          end
          if(_zz_1[3206]) begin
            regVec_3206 <= _zz_regVec_0;
          end
          if(_zz_1[3207]) begin
            regVec_3207 <= _zz_regVec_0;
          end
          if(_zz_1[3208]) begin
            regVec_3208 <= _zz_regVec_0;
          end
          if(_zz_1[3209]) begin
            regVec_3209 <= _zz_regVec_0;
          end
          if(_zz_1[3210]) begin
            regVec_3210 <= _zz_regVec_0;
          end
          if(_zz_1[3211]) begin
            regVec_3211 <= _zz_regVec_0;
          end
          if(_zz_1[3212]) begin
            regVec_3212 <= _zz_regVec_0;
          end
          if(_zz_1[3213]) begin
            regVec_3213 <= _zz_regVec_0;
          end
          if(_zz_1[3214]) begin
            regVec_3214 <= _zz_regVec_0;
          end
          if(_zz_1[3215]) begin
            regVec_3215 <= _zz_regVec_0;
          end
          if(_zz_1[3216]) begin
            regVec_3216 <= _zz_regVec_0;
          end
          if(_zz_1[3217]) begin
            regVec_3217 <= _zz_regVec_0;
          end
          if(_zz_1[3218]) begin
            regVec_3218 <= _zz_regVec_0;
          end
          if(_zz_1[3219]) begin
            regVec_3219 <= _zz_regVec_0;
          end
          if(_zz_1[3220]) begin
            regVec_3220 <= _zz_regVec_0;
          end
          if(_zz_1[3221]) begin
            regVec_3221 <= _zz_regVec_0;
          end
          if(_zz_1[3222]) begin
            regVec_3222 <= _zz_regVec_0;
          end
          if(_zz_1[3223]) begin
            regVec_3223 <= _zz_regVec_0;
          end
          if(_zz_1[3224]) begin
            regVec_3224 <= _zz_regVec_0;
          end
          if(_zz_1[3225]) begin
            regVec_3225 <= _zz_regVec_0;
          end
          if(_zz_1[3226]) begin
            regVec_3226 <= _zz_regVec_0;
          end
          if(_zz_1[3227]) begin
            regVec_3227 <= _zz_regVec_0;
          end
          if(_zz_1[3228]) begin
            regVec_3228 <= _zz_regVec_0;
          end
          if(_zz_1[3229]) begin
            regVec_3229 <= _zz_regVec_0;
          end
          if(_zz_1[3230]) begin
            regVec_3230 <= _zz_regVec_0;
          end
          if(_zz_1[3231]) begin
            regVec_3231 <= _zz_regVec_0;
          end
          if(_zz_1[3232]) begin
            regVec_3232 <= _zz_regVec_0;
          end
          if(_zz_1[3233]) begin
            regVec_3233 <= _zz_regVec_0;
          end
          if(_zz_1[3234]) begin
            regVec_3234 <= _zz_regVec_0;
          end
          if(_zz_1[3235]) begin
            regVec_3235 <= _zz_regVec_0;
          end
          if(_zz_1[3236]) begin
            regVec_3236 <= _zz_regVec_0;
          end
          if(_zz_1[3237]) begin
            regVec_3237 <= _zz_regVec_0;
          end
          if(_zz_1[3238]) begin
            regVec_3238 <= _zz_regVec_0;
          end
          if(_zz_1[3239]) begin
            regVec_3239 <= _zz_regVec_0;
          end
          if(_zz_1[3240]) begin
            regVec_3240 <= _zz_regVec_0;
          end
          if(_zz_1[3241]) begin
            regVec_3241 <= _zz_regVec_0;
          end
          if(_zz_1[3242]) begin
            regVec_3242 <= _zz_regVec_0;
          end
          if(_zz_1[3243]) begin
            regVec_3243 <= _zz_regVec_0;
          end
          if(_zz_1[3244]) begin
            regVec_3244 <= _zz_regVec_0;
          end
          if(_zz_1[3245]) begin
            regVec_3245 <= _zz_regVec_0;
          end
          if(_zz_1[3246]) begin
            regVec_3246 <= _zz_regVec_0;
          end
          if(_zz_1[3247]) begin
            regVec_3247 <= _zz_regVec_0;
          end
          if(_zz_1[3248]) begin
            regVec_3248 <= _zz_regVec_0;
          end
          if(_zz_1[3249]) begin
            regVec_3249 <= _zz_regVec_0;
          end
          if(_zz_1[3250]) begin
            regVec_3250 <= _zz_regVec_0;
          end
          if(_zz_1[3251]) begin
            regVec_3251 <= _zz_regVec_0;
          end
          if(_zz_1[3252]) begin
            regVec_3252 <= _zz_regVec_0;
          end
          if(_zz_1[3253]) begin
            regVec_3253 <= _zz_regVec_0;
          end
          if(_zz_1[3254]) begin
            regVec_3254 <= _zz_regVec_0;
          end
          if(_zz_1[3255]) begin
            regVec_3255 <= _zz_regVec_0;
          end
          if(_zz_1[3256]) begin
            regVec_3256 <= _zz_regVec_0;
          end
          if(_zz_1[3257]) begin
            regVec_3257 <= _zz_regVec_0;
          end
          if(_zz_1[3258]) begin
            regVec_3258 <= _zz_regVec_0;
          end
          if(_zz_1[3259]) begin
            regVec_3259 <= _zz_regVec_0;
          end
          if(_zz_1[3260]) begin
            regVec_3260 <= _zz_regVec_0;
          end
          if(_zz_1[3261]) begin
            regVec_3261 <= _zz_regVec_0;
          end
          if(_zz_1[3262]) begin
            regVec_3262 <= _zz_regVec_0;
          end
          if(_zz_1[3263]) begin
            regVec_3263 <= _zz_regVec_0;
          end
          if(_zz_1[3264]) begin
            regVec_3264 <= _zz_regVec_0;
          end
          if(_zz_1[3265]) begin
            regVec_3265 <= _zz_regVec_0;
          end
          if(_zz_1[3266]) begin
            regVec_3266 <= _zz_regVec_0;
          end
          if(_zz_1[3267]) begin
            regVec_3267 <= _zz_regVec_0;
          end
          if(_zz_1[3268]) begin
            regVec_3268 <= _zz_regVec_0;
          end
          if(_zz_1[3269]) begin
            regVec_3269 <= _zz_regVec_0;
          end
          if(_zz_1[3270]) begin
            regVec_3270 <= _zz_regVec_0;
          end
          if(_zz_1[3271]) begin
            regVec_3271 <= _zz_regVec_0;
          end
          if(_zz_1[3272]) begin
            regVec_3272 <= _zz_regVec_0;
          end
          if(_zz_1[3273]) begin
            regVec_3273 <= _zz_regVec_0;
          end
          if(_zz_1[3274]) begin
            regVec_3274 <= _zz_regVec_0;
          end
          if(_zz_1[3275]) begin
            regVec_3275 <= _zz_regVec_0;
          end
          if(_zz_1[3276]) begin
            regVec_3276 <= _zz_regVec_0;
          end
          if(_zz_1[3277]) begin
            regVec_3277 <= _zz_regVec_0;
          end
          if(_zz_1[3278]) begin
            regVec_3278 <= _zz_regVec_0;
          end
          if(_zz_1[3279]) begin
            regVec_3279 <= _zz_regVec_0;
          end
          if(_zz_1[3280]) begin
            regVec_3280 <= _zz_regVec_0;
          end
          if(_zz_1[3281]) begin
            regVec_3281 <= _zz_regVec_0;
          end
          if(_zz_1[3282]) begin
            regVec_3282 <= _zz_regVec_0;
          end
          if(_zz_1[3283]) begin
            regVec_3283 <= _zz_regVec_0;
          end
          if(_zz_1[3284]) begin
            regVec_3284 <= _zz_regVec_0;
          end
          if(_zz_1[3285]) begin
            regVec_3285 <= _zz_regVec_0;
          end
          if(_zz_1[3286]) begin
            regVec_3286 <= _zz_regVec_0;
          end
          if(_zz_1[3287]) begin
            regVec_3287 <= _zz_regVec_0;
          end
          if(_zz_1[3288]) begin
            regVec_3288 <= _zz_regVec_0;
          end
          if(_zz_1[3289]) begin
            regVec_3289 <= _zz_regVec_0;
          end
          if(_zz_1[3290]) begin
            regVec_3290 <= _zz_regVec_0;
          end
          if(_zz_1[3291]) begin
            regVec_3291 <= _zz_regVec_0;
          end
          if(_zz_1[3292]) begin
            regVec_3292 <= _zz_regVec_0;
          end
          if(_zz_1[3293]) begin
            regVec_3293 <= _zz_regVec_0;
          end
          if(_zz_1[3294]) begin
            regVec_3294 <= _zz_regVec_0;
          end
          if(_zz_1[3295]) begin
            regVec_3295 <= _zz_regVec_0;
          end
          if(_zz_1[3296]) begin
            regVec_3296 <= _zz_regVec_0;
          end
          if(_zz_1[3297]) begin
            regVec_3297 <= _zz_regVec_0;
          end
          if(_zz_1[3298]) begin
            regVec_3298 <= _zz_regVec_0;
          end
          if(_zz_1[3299]) begin
            regVec_3299 <= _zz_regVec_0;
          end
          if(_zz_1[3300]) begin
            regVec_3300 <= _zz_regVec_0;
          end
          if(_zz_1[3301]) begin
            regVec_3301 <= _zz_regVec_0;
          end
          if(_zz_1[3302]) begin
            regVec_3302 <= _zz_regVec_0;
          end
          if(_zz_1[3303]) begin
            regVec_3303 <= _zz_regVec_0;
          end
          if(_zz_1[3304]) begin
            regVec_3304 <= _zz_regVec_0;
          end
          if(_zz_1[3305]) begin
            regVec_3305 <= _zz_regVec_0;
          end
          if(_zz_1[3306]) begin
            regVec_3306 <= _zz_regVec_0;
          end
          if(_zz_1[3307]) begin
            regVec_3307 <= _zz_regVec_0;
          end
          if(_zz_1[3308]) begin
            regVec_3308 <= _zz_regVec_0;
          end
          if(_zz_1[3309]) begin
            regVec_3309 <= _zz_regVec_0;
          end
          if(_zz_1[3310]) begin
            regVec_3310 <= _zz_regVec_0;
          end
          if(_zz_1[3311]) begin
            regVec_3311 <= _zz_regVec_0;
          end
          if(_zz_1[3312]) begin
            regVec_3312 <= _zz_regVec_0;
          end
          if(_zz_1[3313]) begin
            regVec_3313 <= _zz_regVec_0;
          end
          if(_zz_1[3314]) begin
            regVec_3314 <= _zz_regVec_0;
          end
          if(_zz_1[3315]) begin
            regVec_3315 <= _zz_regVec_0;
          end
          if(_zz_1[3316]) begin
            regVec_3316 <= _zz_regVec_0;
          end
          if(_zz_1[3317]) begin
            regVec_3317 <= _zz_regVec_0;
          end
          if(_zz_1[3318]) begin
            regVec_3318 <= _zz_regVec_0;
          end
          if(_zz_1[3319]) begin
            regVec_3319 <= _zz_regVec_0;
          end
          if(_zz_1[3320]) begin
            regVec_3320 <= _zz_regVec_0;
          end
          if(_zz_1[3321]) begin
            regVec_3321 <= _zz_regVec_0;
          end
          if(_zz_1[3322]) begin
            regVec_3322 <= _zz_regVec_0;
          end
          if(_zz_1[3323]) begin
            regVec_3323 <= _zz_regVec_0;
          end
          if(_zz_1[3324]) begin
            regVec_3324 <= _zz_regVec_0;
          end
          if(_zz_1[3325]) begin
            regVec_3325 <= _zz_regVec_0;
          end
          if(_zz_1[3326]) begin
            regVec_3326 <= _zz_regVec_0;
          end
          if(_zz_1[3327]) begin
            regVec_3327 <= _zz_regVec_0;
          end
          if(_zz_1[3328]) begin
            regVec_3328 <= _zz_regVec_0;
          end
          if(_zz_1[3329]) begin
            regVec_3329 <= _zz_regVec_0;
          end
          if(_zz_1[3330]) begin
            regVec_3330 <= _zz_regVec_0;
          end
          if(_zz_1[3331]) begin
            regVec_3331 <= _zz_regVec_0;
          end
          if(_zz_1[3332]) begin
            regVec_3332 <= _zz_regVec_0;
          end
          if(_zz_1[3333]) begin
            regVec_3333 <= _zz_regVec_0;
          end
          if(_zz_1[3334]) begin
            regVec_3334 <= _zz_regVec_0;
          end
          if(_zz_1[3335]) begin
            regVec_3335 <= _zz_regVec_0;
          end
          if(_zz_1[3336]) begin
            regVec_3336 <= _zz_regVec_0;
          end
          if(_zz_1[3337]) begin
            regVec_3337 <= _zz_regVec_0;
          end
          if(_zz_1[3338]) begin
            regVec_3338 <= _zz_regVec_0;
          end
          if(_zz_1[3339]) begin
            regVec_3339 <= _zz_regVec_0;
          end
          if(_zz_1[3340]) begin
            regVec_3340 <= _zz_regVec_0;
          end
          if(_zz_1[3341]) begin
            regVec_3341 <= _zz_regVec_0;
          end
          if(_zz_1[3342]) begin
            regVec_3342 <= _zz_regVec_0;
          end
          if(_zz_1[3343]) begin
            regVec_3343 <= _zz_regVec_0;
          end
          if(_zz_1[3344]) begin
            regVec_3344 <= _zz_regVec_0;
          end
          if(_zz_1[3345]) begin
            regVec_3345 <= _zz_regVec_0;
          end
          if(_zz_1[3346]) begin
            regVec_3346 <= _zz_regVec_0;
          end
          if(_zz_1[3347]) begin
            regVec_3347 <= _zz_regVec_0;
          end
          if(_zz_1[3348]) begin
            regVec_3348 <= _zz_regVec_0;
          end
          if(_zz_1[3349]) begin
            regVec_3349 <= _zz_regVec_0;
          end
          if(_zz_1[3350]) begin
            regVec_3350 <= _zz_regVec_0;
          end
          if(_zz_1[3351]) begin
            regVec_3351 <= _zz_regVec_0;
          end
          if(_zz_1[3352]) begin
            regVec_3352 <= _zz_regVec_0;
          end
          if(_zz_1[3353]) begin
            regVec_3353 <= _zz_regVec_0;
          end
          if(_zz_1[3354]) begin
            regVec_3354 <= _zz_regVec_0;
          end
          if(_zz_1[3355]) begin
            regVec_3355 <= _zz_regVec_0;
          end
          if(_zz_1[3356]) begin
            regVec_3356 <= _zz_regVec_0;
          end
          if(_zz_1[3357]) begin
            regVec_3357 <= _zz_regVec_0;
          end
          if(_zz_1[3358]) begin
            regVec_3358 <= _zz_regVec_0;
          end
          if(_zz_1[3359]) begin
            regVec_3359 <= _zz_regVec_0;
          end
          if(_zz_1[3360]) begin
            regVec_3360 <= _zz_regVec_0;
          end
          if(_zz_1[3361]) begin
            regVec_3361 <= _zz_regVec_0;
          end
          if(_zz_1[3362]) begin
            regVec_3362 <= _zz_regVec_0;
          end
          if(_zz_1[3363]) begin
            regVec_3363 <= _zz_regVec_0;
          end
          if(_zz_1[3364]) begin
            regVec_3364 <= _zz_regVec_0;
          end
          if(_zz_1[3365]) begin
            regVec_3365 <= _zz_regVec_0;
          end
          if(_zz_1[3366]) begin
            regVec_3366 <= _zz_regVec_0;
          end
          if(_zz_1[3367]) begin
            regVec_3367 <= _zz_regVec_0;
          end
          if(_zz_1[3368]) begin
            regVec_3368 <= _zz_regVec_0;
          end
          if(_zz_1[3369]) begin
            regVec_3369 <= _zz_regVec_0;
          end
          if(_zz_1[3370]) begin
            regVec_3370 <= _zz_regVec_0;
          end
          if(_zz_1[3371]) begin
            regVec_3371 <= _zz_regVec_0;
          end
          if(_zz_1[3372]) begin
            regVec_3372 <= _zz_regVec_0;
          end
          if(_zz_1[3373]) begin
            regVec_3373 <= _zz_regVec_0;
          end
          if(_zz_1[3374]) begin
            regVec_3374 <= _zz_regVec_0;
          end
          if(_zz_1[3375]) begin
            regVec_3375 <= _zz_regVec_0;
          end
          if(_zz_1[3376]) begin
            regVec_3376 <= _zz_regVec_0;
          end
          if(_zz_1[3377]) begin
            regVec_3377 <= _zz_regVec_0;
          end
          if(_zz_1[3378]) begin
            regVec_3378 <= _zz_regVec_0;
          end
          if(_zz_1[3379]) begin
            regVec_3379 <= _zz_regVec_0;
          end
          if(_zz_1[3380]) begin
            regVec_3380 <= _zz_regVec_0;
          end
          if(_zz_1[3381]) begin
            regVec_3381 <= _zz_regVec_0;
          end
          if(_zz_1[3382]) begin
            regVec_3382 <= _zz_regVec_0;
          end
          if(_zz_1[3383]) begin
            regVec_3383 <= _zz_regVec_0;
          end
          if(_zz_1[3384]) begin
            regVec_3384 <= _zz_regVec_0;
          end
          if(_zz_1[3385]) begin
            regVec_3385 <= _zz_regVec_0;
          end
          if(_zz_1[3386]) begin
            regVec_3386 <= _zz_regVec_0;
          end
          if(_zz_1[3387]) begin
            regVec_3387 <= _zz_regVec_0;
          end
          if(_zz_1[3388]) begin
            regVec_3388 <= _zz_regVec_0;
          end
          if(_zz_1[3389]) begin
            regVec_3389 <= _zz_regVec_0;
          end
          if(_zz_1[3390]) begin
            regVec_3390 <= _zz_regVec_0;
          end
          if(_zz_1[3391]) begin
            regVec_3391 <= _zz_regVec_0;
          end
          if(_zz_1[3392]) begin
            regVec_3392 <= _zz_regVec_0;
          end
          if(_zz_1[3393]) begin
            regVec_3393 <= _zz_regVec_0;
          end
          if(_zz_1[3394]) begin
            regVec_3394 <= _zz_regVec_0;
          end
          if(_zz_1[3395]) begin
            regVec_3395 <= _zz_regVec_0;
          end
          if(_zz_1[3396]) begin
            regVec_3396 <= _zz_regVec_0;
          end
          if(_zz_1[3397]) begin
            regVec_3397 <= _zz_regVec_0;
          end
          if(_zz_1[3398]) begin
            regVec_3398 <= _zz_regVec_0;
          end
          if(_zz_1[3399]) begin
            regVec_3399 <= _zz_regVec_0;
          end
          if(_zz_1[3400]) begin
            regVec_3400 <= _zz_regVec_0;
          end
          if(_zz_1[3401]) begin
            regVec_3401 <= _zz_regVec_0;
          end
          if(_zz_1[3402]) begin
            regVec_3402 <= _zz_regVec_0;
          end
          if(_zz_1[3403]) begin
            regVec_3403 <= _zz_regVec_0;
          end
          if(_zz_1[3404]) begin
            regVec_3404 <= _zz_regVec_0;
          end
          if(_zz_1[3405]) begin
            regVec_3405 <= _zz_regVec_0;
          end
          if(_zz_1[3406]) begin
            regVec_3406 <= _zz_regVec_0;
          end
          if(_zz_1[3407]) begin
            regVec_3407 <= _zz_regVec_0;
          end
          if(_zz_1[3408]) begin
            regVec_3408 <= _zz_regVec_0;
          end
          if(_zz_1[3409]) begin
            regVec_3409 <= _zz_regVec_0;
          end
          if(_zz_1[3410]) begin
            regVec_3410 <= _zz_regVec_0;
          end
          if(_zz_1[3411]) begin
            regVec_3411 <= _zz_regVec_0;
          end
          if(_zz_1[3412]) begin
            regVec_3412 <= _zz_regVec_0;
          end
          if(_zz_1[3413]) begin
            regVec_3413 <= _zz_regVec_0;
          end
          if(_zz_1[3414]) begin
            regVec_3414 <= _zz_regVec_0;
          end
          if(_zz_1[3415]) begin
            regVec_3415 <= _zz_regVec_0;
          end
          if(_zz_1[3416]) begin
            regVec_3416 <= _zz_regVec_0;
          end
          if(_zz_1[3417]) begin
            regVec_3417 <= _zz_regVec_0;
          end
          if(_zz_1[3418]) begin
            regVec_3418 <= _zz_regVec_0;
          end
          if(_zz_1[3419]) begin
            regVec_3419 <= _zz_regVec_0;
          end
          if(_zz_1[3420]) begin
            regVec_3420 <= _zz_regVec_0;
          end
          if(_zz_1[3421]) begin
            regVec_3421 <= _zz_regVec_0;
          end
          if(_zz_1[3422]) begin
            regVec_3422 <= _zz_regVec_0;
          end
          if(_zz_1[3423]) begin
            regVec_3423 <= _zz_regVec_0;
          end
          if(_zz_1[3424]) begin
            regVec_3424 <= _zz_regVec_0;
          end
          if(_zz_1[3425]) begin
            regVec_3425 <= _zz_regVec_0;
          end
          if(_zz_1[3426]) begin
            regVec_3426 <= _zz_regVec_0;
          end
          if(_zz_1[3427]) begin
            regVec_3427 <= _zz_regVec_0;
          end
          if(_zz_1[3428]) begin
            regVec_3428 <= _zz_regVec_0;
          end
          if(_zz_1[3429]) begin
            regVec_3429 <= _zz_regVec_0;
          end
          if(_zz_1[3430]) begin
            regVec_3430 <= _zz_regVec_0;
          end
          if(_zz_1[3431]) begin
            regVec_3431 <= _zz_regVec_0;
          end
          if(_zz_1[3432]) begin
            regVec_3432 <= _zz_regVec_0;
          end
          if(_zz_1[3433]) begin
            regVec_3433 <= _zz_regVec_0;
          end
          if(_zz_1[3434]) begin
            regVec_3434 <= _zz_regVec_0;
          end
          if(_zz_1[3435]) begin
            regVec_3435 <= _zz_regVec_0;
          end
          if(_zz_1[3436]) begin
            regVec_3436 <= _zz_regVec_0;
          end
          if(_zz_1[3437]) begin
            regVec_3437 <= _zz_regVec_0;
          end
          if(_zz_1[3438]) begin
            regVec_3438 <= _zz_regVec_0;
          end
          if(_zz_1[3439]) begin
            regVec_3439 <= _zz_regVec_0;
          end
          if(_zz_1[3440]) begin
            regVec_3440 <= _zz_regVec_0;
          end
          if(_zz_1[3441]) begin
            regVec_3441 <= _zz_regVec_0;
          end
          if(_zz_1[3442]) begin
            regVec_3442 <= _zz_regVec_0;
          end
          if(_zz_1[3443]) begin
            regVec_3443 <= _zz_regVec_0;
          end
          if(_zz_1[3444]) begin
            regVec_3444 <= _zz_regVec_0;
          end
          if(_zz_1[3445]) begin
            regVec_3445 <= _zz_regVec_0;
          end
          if(_zz_1[3446]) begin
            regVec_3446 <= _zz_regVec_0;
          end
          if(_zz_1[3447]) begin
            regVec_3447 <= _zz_regVec_0;
          end
          if(_zz_1[3448]) begin
            regVec_3448 <= _zz_regVec_0;
          end
          if(_zz_1[3449]) begin
            regVec_3449 <= _zz_regVec_0;
          end
          if(_zz_1[3450]) begin
            regVec_3450 <= _zz_regVec_0;
          end
          if(_zz_1[3451]) begin
            regVec_3451 <= _zz_regVec_0;
          end
          if(_zz_1[3452]) begin
            regVec_3452 <= _zz_regVec_0;
          end
          if(_zz_1[3453]) begin
            regVec_3453 <= _zz_regVec_0;
          end
          if(_zz_1[3454]) begin
            regVec_3454 <= _zz_regVec_0;
          end
          if(_zz_1[3455]) begin
            regVec_3455 <= _zz_regVec_0;
          end
          if(_zz_1[3456]) begin
            regVec_3456 <= _zz_regVec_0;
          end
          if(_zz_1[3457]) begin
            regVec_3457 <= _zz_regVec_0;
          end
          if(_zz_1[3458]) begin
            regVec_3458 <= _zz_regVec_0;
          end
          if(_zz_1[3459]) begin
            regVec_3459 <= _zz_regVec_0;
          end
          if(_zz_1[3460]) begin
            regVec_3460 <= _zz_regVec_0;
          end
          if(_zz_1[3461]) begin
            regVec_3461 <= _zz_regVec_0;
          end
          if(_zz_1[3462]) begin
            regVec_3462 <= _zz_regVec_0;
          end
          if(_zz_1[3463]) begin
            regVec_3463 <= _zz_regVec_0;
          end
          if(_zz_1[3464]) begin
            regVec_3464 <= _zz_regVec_0;
          end
          if(_zz_1[3465]) begin
            regVec_3465 <= _zz_regVec_0;
          end
          if(_zz_1[3466]) begin
            regVec_3466 <= _zz_regVec_0;
          end
          if(_zz_1[3467]) begin
            regVec_3467 <= _zz_regVec_0;
          end
          if(_zz_1[3468]) begin
            regVec_3468 <= _zz_regVec_0;
          end
          if(_zz_1[3469]) begin
            regVec_3469 <= _zz_regVec_0;
          end
          if(_zz_1[3470]) begin
            regVec_3470 <= _zz_regVec_0;
          end
          if(_zz_1[3471]) begin
            regVec_3471 <= _zz_regVec_0;
          end
          if(_zz_1[3472]) begin
            regVec_3472 <= _zz_regVec_0;
          end
          if(_zz_1[3473]) begin
            regVec_3473 <= _zz_regVec_0;
          end
          if(_zz_1[3474]) begin
            regVec_3474 <= _zz_regVec_0;
          end
          if(_zz_1[3475]) begin
            regVec_3475 <= _zz_regVec_0;
          end
          if(_zz_1[3476]) begin
            regVec_3476 <= _zz_regVec_0;
          end
          if(_zz_1[3477]) begin
            regVec_3477 <= _zz_regVec_0;
          end
          if(_zz_1[3478]) begin
            regVec_3478 <= _zz_regVec_0;
          end
          if(_zz_1[3479]) begin
            regVec_3479 <= _zz_regVec_0;
          end
          if(_zz_1[3480]) begin
            regVec_3480 <= _zz_regVec_0;
          end
          if(_zz_1[3481]) begin
            regVec_3481 <= _zz_regVec_0;
          end
          if(_zz_1[3482]) begin
            regVec_3482 <= _zz_regVec_0;
          end
          if(_zz_1[3483]) begin
            regVec_3483 <= _zz_regVec_0;
          end
          if(_zz_1[3484]) begin
            regVec_3484 <= _zz_regVec_0;
          end
          if(_zz_1[3485]) begin
            regVec_3485 <= _zz_regVec_0;
          end
          if(_zz_1[3486]) begin
            regVec_3486 <= _zz_regVec_0;
          end
          if(_zz_1[3487]) begin
            regVec_3487 <= _zz_regVec_0;
          end
          if(_zz_1[3488]) begin
            regVec_3488 <= _zz_regVec_0;
          end
          if(_zz_1[3489]) begin
            regVec_3489 <= _zz_regVec_0;
          end
          if(_zz_1[3490]) begin
            regVec_3490 <= _zz_regVec_0;
          end
          if(_zz_1[3491]) begin
            regVec_3491 <= _zz_regVec_0;
          end
          if(_zz_1[3492]) begin
            regVec_3492 <= _zz_regVec_0;
          end
          if(_zz_1[3493]) begin
            regVec_3493 <= _zz_regVec_0;
          end
          if(_zz_1[3494]) begin
            regVec_3494 <= _zz_regVec_0;
          end
          if(_zz_1[3495]) begin
            regVec_3495 <= _zz_regVec_0;
          end
          if(_zz_1[3496]) begin
            regVec_3496 <= _zz_regVec_0;
          end
          if(_zz_1[3497]) begin
            regVec_3497 <= _zz_regVec_0;
          end
          if(_zz_1[3498]) begin
            regVec_3498 <= _zz_regVec_0;
          end
          if(_zz_1[3499]) begin
            regVec_3499 <= _zz_regVec_0;
          end
          if(_zz_1[3500]) begin
            regVec_3500 <= _zz_regVec_0;
          end
          if(_zz_1[3501]) begin
            regVec_3501 <= _zz_regVec_0;
          end
          if(_zz_1[3502]) begin
            regVec_3502 <= _zz_regVec_0;
          end
          if(_zz_1[3503]) begin
            regVec_3503 <= _zz_regVec_0;
          end
          if(_zz_1[3504]) begin
            regVec_3504 <= _zz_regVec_0;
          end
          if(_zz_1[3505]) begin
            regVec_3505 <= _zz_regVec_0;
          end
          if(_zz_1[3506]) begin
            regVec_3506 <= _zz_regVec_0;
          end
          if(_zz_1[3507]) begin
            regVec_3507 <= _zz_regVec_0;
          end
          if(_zz_1[3508]) begin
            regVec_3508 <= _zz_regVec_0;
          end
          if(_zz_1[3509]) begin
            regVec_3509 <= _zz_regVec_0;
          end
          if(_zz_1[3510]) begin
            regVec_3510 <= _zz_regVec_0;
          end
          if(_zz_1[3511]) begin
            regVec_3511 <= _zz_regVec_0;
          end
          if(_zz_1[3512]) begin
            regVec_3512 <= _zz_regVec_0;
          end
          if(_zz_1[3513]) begin
            regVec_3513 <= _zz_regVec_0;
          end
          if(_zz_1[3514]) begin
            regVec_3514 <= _zz_regVec_0;
          end
          if(_zz_1[3515]) begin
            regVec_3515 <= _zz_regVec_0;
          end
          if(_zz_1[3516]) begin
            regVec_3516 <= _zz_regVec_0;
          end
          if(_zz_1[3517]) begin
            regVec_3517 <= _zz_regVec_0;
          end
          if(_zz_1[3518]) begin
            regVec_3518 <= _zz_regVec_0;
          end
          if(_zz_1[3519]) begin
            regVec_3519 <= _zz_regVec_0;
          end
          if(_zz_1[3520]) begin
            regVec_3520 <= _zz_regVec_0;
          end
          if(_zz_1[3521]) begin
            regVec_3521 <= _zz_regVec_0;
          end
          if(_zz_1[3522]) begin
            regVec_3522 <= _zz_regVec_0;
          end
          if(_zz_1[3523]) begin
            regVec_3523 <= _zz_regVec_0;
          end
          if(_zz_1[3524]) begin
            regVec_3524 <= _zz_regVec_0;
          end
          if(_zz_1[3525]) begin
            regVec_3525 <= _zz_regVec_0;
          end
          if(_zz_1[3526]) begin
            regVec_3526 <= _zz_regVec_0;
          end
          if(_zz_1[3527]) begin
            regVec_3527 <= _zz_regVec_0;
          end
          if(_zz_1[3528]) begin
            regVec_3528 <= _zz_regVec_0;
          end
          if(_zz_1[3529]) begin
            regVec_3529 <= _zz_regVec_0;
          end
          if(_zz_1[3530]) begin
            regVec_3530 <= _zz_regVec_0;
          end
          if(_zz_1[3531]) begin
            regVec_3531 <= _zz_regVec_0;
          end
          if(_zz_1[3532]) begin
            regVec_3532 <= _zz_regVec_0;
          end
          if(_zz_1[3533]) begin
            regVec_3533 <= _zz_regVec_0;
          end
          if(_zz_1[3534]) begin
            regVec_3534 <= _zz_regVec_0;
          end
          if(_zz_1[3535]) begin
            regVec_3535 <= _zz_regVec_0;
          end
          if(_zz_1[3536]) begin
            regVec_3536 <= _zz_regVec_0;
          end
          if(_zz_1[3537]) begin
            regVec_3537 <= _zz_regVec_0;
          end
          if(_zz_1[3538]) begin
            regVec_3538 <= _zz_regVec_0;
          end
          if(_zz_1[3539]) begin
            regVec_3539 <= _zz_regVec_0;
          end
          if(_zz_1[3540]) begin
            regVec_3540 <= _zz_regVec_0;
          end
          if(_zz_1[3541]) begin
            regVec_3541 <= _zz_regVec_0;
          end
          if(_zz_1[3542]) begin
            regVec_3542 <= _zz_regVec_0;
          end
          if(_zz_1[3543]) begin
            regVec_3543 <= _zz_regVec_0;
          end
          if(_zz_1[3544]) begin
            regVec_3544 <= _zz_regVec_0;
          end
          if(_zz_1[3545]) begin
            regVec_3545 <= _zz_regVec_0;
          end
          if(_zz_1[3546]) begin
            regVec_3546 <= _zz_regVec_0;
          end
          if(_zz_1[3547]) begin
            regVec_3547 <= _zz_regVec_0;
          end
          if(_zz_1[3548]) begin
            regVec_3548 <= _zz_regVec_0;
          end
          if(_zz_1[3549]) begin
            regVec_3549 <= _zz_regVec_0;
          end
          if(_zz_1[3550]) begin
            regVec_3550 <= _zz_regVec_0;
          end
          if(_zz_1[3551]) begin
            regVec_3551 <= _zz_regVec_0;
          end
          if(_zz_1[3552]) begin
            regVec_3552 <= _zz_regVec_0;
          end
          if(_zz_1[3553]) begin
            regVec_3553 <= _zz_regVec_0;
          end
          if(_zz_1[3554]) begin
            regVec_3554 <= _zz_regVec_0;
          end
          if(_zz_1[3555]) begin
            regVec_3555 <= _zz_regVec_0;
          end
          if(_zz_1[3556]) begin
            regVec_3556 <= _zz_regVec_0;
          end
          if(_zz_1[3557]) begin
            regVec_3557 <= _zz_regVec_0;
          end
          if(_zz_1[3558]) begin
            regVec_3558 <= _zz_regVec_0;
          end
          if(_zz_1[3559]) begin
            regVec_3559 <= _zz_regVec_0;
          end
          if(_zz_1[3560]) begin
            regVec_3560 <= _zz_regVec_0;
          end
          if(_zz_1[3561]) begin
            regVec_3561 <= _zz_regVec_0;
          end
          if(_zz_1[3562]) begin
            regVec_3562 <= _zz_regVec_0;
          end
          if(_zz_1[3563]) begin
            regVec_3563 <= _zz_regVec_0;
          end
          if(_zz_1[3564]) begin
            regVec_3564 <= _zz_regVec_0;
          end
          if(_zz_1[3565]) begin
            regVec_3565 <= _zz_regVec_0;
          end
          if(_zz_1[3566]) begin
            regVec_3566 <= _zz_regVec_0;
          end
          if(_zz_1[3567]) begin
            regVec_3567 <= _zz_regVec_0;
          end
          if(_zz_1[3568]) begin
            regVec_3568 <= _zz_regVec_0;
          end
          if(_zz_1[3569]) begin
            regVec_3569 <= _zz_regVec_0;
          end
          if(_zz_1[3570]) begin
            regVec_3570 <= _zz_regVec_0;
          end
          if(_zz_1[3571]) begin
            regVec_3571 <= _zz_regVec_0;
          end
          if(_zz_1[3572]) begin
            regVec_3572 <= _zz_regVec_0;
          end
          if(_zz_1[3573]) begin
            regVec_3573 <= _zz_regVec_0;
          end
          if(_zz_1[3574]) begin
            regVec_3574 <= _zz_regVec_0;
          end
          if(_zz_1[3575]) begin
            regVec_3575 <= _zz_regVec_0;
          end
          if(_zz_1[3576]) begin
            regVec_3576 <= _zz_regVec_0;
          end
          if(_zz_1[3577]) begin
            regVec_3577 <= _zz_regVec_0;
          end
          if(_zz_1[3578]) begin
            regVec_3578 <= _zz_regVec_0;
          end
          if(_zz_1[3579]) begin
            regVec_3579 <= _zz_regVec_0;
          end
          if(_zz_1[3580]) begin
            regVec_3580 <= _zz_regVec_0;
          end
          if(_zz_1[3581]) begin
            regVec_3581 <= _zz_regVec_0;
          end
          if(_zz_1[3582]) begin
            regVec_3582 <= _zz_regVec_0;
          end
          if(_zz_1[3583]) begin
            regVec_3583 <= _zz_regVec_0;
          end
          if(_zz_1[3584]) begin
            regVec_3584 <= _zz_regVec_0;
          end
          if(_zz_1[3585]) begin
            regVec_3585 <= _zz_regVec_0;
          end
          if(_zz_1[3586]) begin
            regVec_3586 <= _zz_regVec_0;
          end
          if(_zz_1[3587]) begin
            regVec_3587 <= _zz_regVec_0;
          end
          if(_zz_1[3588]) begin
            regVec_3588 <= _zz_regVec_0;
          end
          if(_zz_1[3589]) begin
            regVec_3589 <= _zz_regVec_0;
          end
          if(_zz_1[3590]) begin
            regVec_3590 <= _zz_regVec_0;
          end
          if(_zz_1[3591]) begin
            regVec_3591 <= _zz_regVec_0;
          end
          if(_zz_1[3592]) begin
            regVec_3592 <= _zz_regVec_0;
          end
          if(_zz_1[3593]) begin
            regVec_3593 <= _zz_regVec_0;
          end
          if(_zz_1[3594]) begin
            regVec_3594 <= _zz_regVec_0;
          end
          if(_zz_1[3595]) begin
            regVec_3595 <= _zz_regVec_0;
          end
          if(_zz_1[3596]) begin
            regVec_3596 <= _zz_regVec_0;
          end
          if(_zz_1[3597]) begin
            regVec_3597 <= _zz_regVec_0;
          end
          if(_zz_1[3598]) begin
            regVec_3598 <= _zz_regVec_0;
          end
          if(_zz_1[3599]) begin
            regVec_3599 <= _zz_regVec_0;
          end
          if(_zz_1[3600]) begin
            regVec_3600 <= _zz_regVec_0;
          end
          if(_zz_1[3601]) begin
            regVec_3601 <= _zz_regVec_0;
          end
          if(_zz_1[3602]) begin
            regVec_3602 <= _zz_regVec_0;
          end
          if(_zz_1[3603]) begin
            regVec_3603 <= _zz_regVec_0;
          end
          if(_zz_1[3604]) begin
            regVec_3604 <= _zz_regVec_0;
          end
          if(_zz_1[3605]) begin
            regVec_3605 <= _zz_regVec_0;
          end
          if(_zz_1[3606]) begin
            regVec_3606 <= _zz_regVec_0;
          end
          if(_zz_1[3607]) begin
            regVec_3607 <= _zz_regVec_0;
          end
          if(_zz_1[3608]) begin
            regVec_3608 <= _zz_regVec_0;
          end
          if(_zz_1[3609]) begin
            regVec_3609 <= _zz_regVec_0;
          end
          if(_zz_1[3610]) begin
            regVec_3610 <= _zz_regVec_0;
          end
          if(_zz_1[3611]) begin
            regVec_3611 <= _zz_regVec_0;
          end
          if(_zz_1[3612]) begin
            regVec_3612 <= _zz_regVec_0;
          end
          if(_zz_1[3613]) begin
            regVec_3613 <= _zz_regVec_0;
          end
          if(_zz_1[3614]) begin
            regVec_3614 <= _zz_regVec_0;
          end
          if(_zz_1[3615]) begin
            regVec_3615 <= _zz_regVec_0;
          end
          if(_zz_1[3616]) begin
            regVec_3616 <= _zz_regVec_0;
          end
          if(_zz_1[3617]) begin
            regVec_3617 <= _zz_regVec_0;
          end
          if(_zz_1[3618]) begin
            regVec_3618 <= _zz_regVec_0;
          end
          if(_zz_1[3619]) begin
            regVec_3619 <= _zz_regVec_0;
          end
          if(_zz_1[3620]) begin
            regVec_3620 <= _zz_regVec_0;
          end
          if(_zz_1[3621]) begin
            regVec_3621 <= _zz_regVec_0;
          end
          if(_zz_1[3622]) begin
            regVec_3622 <= _zz_regVec_0;
          end
          if(_zz_1[3623]) begin
            regVec_3623 <= _zz_regVec_0;
          end
          if(_zz_1[3624]) begin
            regVec_3624 <= _zz_regVec_0;
          end
          if(_zz_1[3625]) begin
            regVec_3625 <= _zz_regVec_0;
          end
          if(_zz_1[3626]) begin
            regVec_3626 <= _zz_regVec_0;
          end
          if(_zz_1[3627]) begin
            regVec_3627 <= _zz_regVec_0;
          end
          if(_zz_1[3628]) begin
            regVec_3628 <= _zz_regVec_0;
          end
          if(_zz_1[3629]) begin
            regVec_3629 <= _zz_regVec_0;
          end
          if(_zz_1[3630]) begin
            regVec_3630 <= _zz_regVec_0;
          end
          if(_zz_1[3631]) begin
            regVec_3631 <= _zz_regVec_0;
          end
          if(_zz_1[3632]) begin
            regVec_3632 <= _zz_regVec_0;
          end
          if(_zz_1[3633]) begin
            regVec_3633 <= _zz_regVec_0;
          end
          if(_zz_1[3634]) begin
            regVec_3634 <= _zz_regVec_0;
          end
          if(_zz_1[3635]) begin
            regVec_3635 <= _zz_regVec_0;
          end
          if(_zz_1[3636]) begin
            regVec_3636 <= _zz_regVec_0;
          end
          if(_zz_1[3637]) begin
            regVec_3637 <= _zz_regVec_0;
          end
          if(_zz_1[3638]) begin
            regVec_3638 <= _zz_regVec_0;
          end
          if(_zz_1[3639]) begin
            regVec_3639 <= _zz_regVec_0;
          end
          if(_zz_1[3640]) begin
            regVec_3640 <= _zz_regVec_0;
          end
          if(_zz_1[3641]) begin
            regVec_3641 <= _zz_regVec_0;
          end
          if(_zz_1[3642]) begin
            regVec_3642 <= _zz_regVec_0;
          end
          if(_zz_1[3643]) begin
            regVec_3643 <= _zz_regVec_0;
          end
          if(_zz_1[3644]) begin
            regVec_3644 <= _zz_regVec_0;
          end
          if(_zz_1[3645]) begin
            regVec_3645 <= _zz_regVec_0;
          end
          if(_zz_1[3646]) begin
            regVec_3646 <= _zz_regVec_0;
          end
          if(_zz_1[3647]) begin
            regVec_3647 <= _zz_regVec_0;
          end
          if(_zz_1[3648]) begin
            regVec_3648 <= _zz_regVec_0;
          end
          if(_zz_1[3649]) begin
            regVec_3649 <= _zz_regVec_0;
          end
          if(_zz_1[3650]) begin
            regVec_3650 <= _zz_regVec_0;
          end
          if(_zz_1[3651]) begin
            regVec_3651 <= _zz_regVec_0;
          end
          if(_zz_1[3652]) begin
            regVec_3652 <= _zz_regVec_0;
          end
          if(_zz_1[3653]) begin
            regVec_3653 <= _zz_regVec_0;
          end
          if(_zz_1[3654]) begin
            regVec_3654 <= _zz_regVec_0;
          end
          if(_zz_1[3655]) begin
            regVec_3655 <= _zz_regVec_0;
          end
          if(_zz_1[3656]) begin
            regVec_3656 <= _zz_regVec_0;
          end
          if(_zz_1[3657]) begin
            regVec_3657 <= _zz_regVec_0;
          end
          if(_zz_1[3658]) begin
            regVec_3658 <= _zz_regVec_0;
          end
          if(_zz_1[3659]) begin
            regVec_3659 <= _zz_regVec_0;
          end
          if(_zz_1[3660]) begin
            regVec_3660 <= _zz_regVec_0;
          end
          if(_zz_1[3661]) begin
            regVec_3661 <= _zz_regVec_0;
          end
          if(_zz_1[3662]) begin
            regVec_3662 <= _zz_regVec_0;
          end
          if(_zz_1[3663]) begin
            regVec_3663 <= _zz_regVec_0;
          end
          if(_zz_1[3664]) begin
            regVec_3664 <= _zz_regVec_0;
          end
          if(_zz_1[3665]) begin
            regVec_3665 <= _zz_regVec_0;
          end
          if(_zz_1[3666]) begin
            regVec_3666 <= _zz_regVec_0;
          end
          if(_zz_1[3667]) begin
            regVec_3667 <= _zz_regVec_0;
          end
          if(_zz_1[3668]) begin
            regVec_3668 <= _zz_regVec_0;
          end
          if(_zz_1[3669]) begin
            regVec_3669 <= _zz_regVec_0;
          end
          if(_zz_1[3670]) begin
            regVec_3670 <= _zz_regVec_0;
          end
          if(_zz_1[3671]) begin
            regVec_3671 <= _zz_regVec_0;
          end
          if(_zz_1[3672]) begin
            regVec_3672 <= _zz_regVec_0;
          end
          if(_zz_1[3673]) begin
            regVec_3673 <= _zz_regVec_0;
          end
          if(_zz_1[3674]) begin
            regVec_3674 <= _zz_regVec_0;
          end
          if(_zz_1[3675]) begin
            regVec_3675 <= _zz_regVec_0;
          end
          if(_zz_1[3676]) begin
            regVec_3676 <= _zz_regVec_0;
          end
          if(_zz_1[3677]) begin
            regVec_3677 <= _zz_regVec_0;
          end
          if(_zz_1[3678]) begin
            regVec_3678 <= _zz_regVec_0;
          end
          if(_zz_1[3679]) begin
            regVec_3679 <= _zz_regVec_0;
          end
          if(_zz_1[3680]) begin
            regVec_3680 <= _zz_regVec_0;
          end
          if(_zz_1[3681]) begin
            regVec_3681 <= _zz_regVec_0;
          end
          if(_zz_1[3682]) begin
            regVec_3682 <= _zz_regVec_0;
          end
          if(_zz_1[3683]) begin
            regVec_3683 <= _zz_regVec_0;
          end
          if(_zz_1[3684]) begin
            regVec_3684 <= _zz_regVec_0;
          end
          if(_zz_1[3685]) begin
            regVec_3685 <= _zz_regVec_0;
          end
          if(_zz_1[3686]) begin
            regVec_3686 <= _zz_regVec_0;
          end
          if(_zz_1[3687]) begin
            regVec_3687 <= _zz_regVec_0;
          end
          if(_zz_1[3688]) begin
            regVec_3688 <= _zz_regVec_0;
          end
          if(_zz_1[3689]) begin
            regVec_3689 <= _zz_regVec_0;
          end
          if(_zz_1[3690]) begin
            regVec_3690 <= _zz_regVec_0;
          end
          if(_zz_1[3691]) begin
            regVec_3691 <= _zz_regVec_0;
          end
          if(_zz_1[3692]) begin
            regVec_3692 <= _zz_regVec_0;
          end
          if(_zz_1[3693]) begin
            regVec_3693 <= _zz_regVec_0;
          end
          if(_zz_1[3694]) begin
            regVec_3694 <= _zz_regVec_0;
          end
          if(_zz_1[3695]) begin
            regVec_3695 <= _zz_regVec_0;
          end
          if(_zz_1[3696]) begin
            regVec_3696 <= _zz_regVec_0;
          end
          if(_zz_1[3697]) begin
            regVec_3697 <= _zz_regVec_0;
          end
          if(_zz_1[3698]) begin
            regVec_3698 <= _zz_regVec_0;
          end
          if(_zz_1[3699]) begin
            regVec_3699 <= _zz_regVec_0;
          end
          if(_zz_1[3700]) begin
            regVec_3700 <= _zz_regVec_0;
          end
          if(_zz_1[3701]) begin
            regVec_3701 <= _zz_regVec_0;
          end
          if(_zz_1[3702]) begin
            regVec_3702 <= _zz_regVec_0;
          end
          if(_zz_1[3703]) begin
            regVec_3703 <= _zz_regVec_0;
          end
          if(_zz_1[3704]) begin
            regVec_3704 <= _zz_regVec_0;
          end
          if(_zz_1[3705]) begin
            regVec_3705 <= _zz_regVec_0;
          end
          if(_zz_1[3706]) begin
            regVec_3706 <= _zz_regVec_0;
          end
          if(_zz_1[3707]) begin
            regVec_3707 <= _zz_regVec_0;
          end
          if(_zz_1[3708]) begin
            regVec_3708 <= _zz_regVec_0;
          end
          if(_zz_1[3709]) begin
            regVec_3709 <= _zz_regVec_0;
          end
          if(_zz_1[3710]) begin
            regVec_3710 <= _zz_regVec_0;
          end
          if(_zz_1[3711]) begin
            regVec_3711 <= _zz_regVec_0;
          end
          if(_zz_1[3712]) begin
            regVec_3712 <= _zz_regVec_0;
          end
          if(_zz_1[3713]) begin
            regVec_3713 <= _zz_regVec_0;
          end
          if(_zz_1[3714]) begin
            regVec_3714 <= _zz_regVec_0;
          end
          if(_zz_1[3715]) begin
            regVec_3715 <= _zz_regVec_0;
          end
          if(_zz_1[3716]) begin
            regVec_3716 <= _zz_regVec_0;
          end
          if(_zz_1[3717]) begin
            regVec_3717 <= _zz_regVec_0;
          end
          if(_zz_1[3718]) begin
            regVec_3718 <= _zz_regVec_0;
          end
          if(_zz_1[3719]) begin
            regVec_3719 <= _zz_regVec_0;
          end
          if(_zz_1[3720]) begin
            regVec_3720 <= _zz_regVec_0;
          end
          if(_zz_1[3721]) begin
            regVec_3721 <= _zz_regVec_0;
          end
          if(_zz_1[3722]) begin
            regVec_3722 <= _zz_regVec_0;
          end
          if(_zz_1[3723]) begin
            regVec_3723 <= _zz_regVec_0;
          end
          if(_zz_1[3724]) begin
            regVec_3724 <= _zz_regVec_0;
          end
          if(_zz_1[3725]) begin
            regVec_3725 <= _zz_regVec_0;
          end
          if(_zz_1[3726]) begin
            regVec_3726 <= _zz_regVec_0;
          end
          if(_zz_1[3727]) begin
            regVec_3727 <= _zz_regVec_0;
          end
          if(_zz_1[3728]) begin
            regVec_3728 <= _zz_regVec_0;
          end
          if(_zz_1[3729]) begin
            regVec_3729 <= _zz_regVec_0;
          end
          if(_zz_1[3730]) begin
            regVec_3730 <= _zz_regVec_0;
          end
          if(_zz_1[3731]) begin
            regVec_3731 <= _zz_regVec_0;
          end
          if(_zz_1[3732]) begin
            regVec_3732 <= _zz_regVec_0;
          end
          if(_zz_1[3733]) begin
            regVec_3733 <= _zz_regVec_0;
          end
          if(_zz_1[3734]) begin
            regVec_3734 <= _zz_regVec_0;
          end
          if(_zz_1[3735]) begin
            regVec_3735 <= _zz_regVec_0;
          end
          if(_zz_1[3736]) begin
            regVec_3736 <= _zz_regVec_0;
          end
          if(_zz_1[3737]) begin
            regVec_3737 <= _zz_regVec_0;
          end
          if(_zz_1[3738]) begin
            regVec_3738 <= _zz_regVec_0;
          end
          if(_zz_1[3739]) begin
            regVec_3739 <= _zz_regVec_0;
          end
          if(_zz_1[3740]) begin
            regVec_3740 <= _zz_regVec_0;
          end
          if(_zz_1[3741]) begin
            regVec_3741 <= _zz_regVec_0;
          end
          if(_zz_1[3742]) begin
            regVec_3742 <= _zz_regVec_0;
          end
          if(_zz_1[3743]) begin
            regVec_3743 <= _zz_regVec_0;
          end
          if(_zz_1[3744]) begin
            regVec_3744 <= _zz_regVec_0;
          end
          if(_zz_1[3745]) begin
            regVec_3745 <= _zz_regVec_0;
          end
          if(_zz_1[3746]) begin
            regVec_3746 <= _zz_regVec_0;
          end
          if(_zz_1[3747]) begin
            regVec_3747 <= _zz_regVec_0;
          end
          if(_zz_1[3748]) begin
            regVec_3748 <= _zz_regVec_0;
          end
          if(_zz_1[3749]) begin
            regVec_3749 <= _zz_regVec_0;
          end
          if(_zz_1[3750]) begin
            regVec_3750 <= _zz_regVec_0;
          end
          if(_zz_1[3751]) begin
            regVec_3751 <= _zz_regVec_0;
          end
          if(_zz_1[3752]) begin
            regVec_3752 <= _zz_regVec_0;
          end
          if(_zz_1[3753]) begin
            regVec_3753 <= _zz_regVec_0;
          end
          if(_zz_1[3754]) begin
            regVec_3754 <= _zz_regVec_0;
          end
          if(_zz_1[3755]) begin
            regVec_3755 <= _zz_regVec_0;
          end
          if(_zz_1[3756]) begin
            regVec_3756 <= _zz_regVec_0;
          end
          if(_zz_1[3757]) begin
            regVec_3757 <= _zz_regVec_0;
          end
          if(_zz_1[3758]) begin
            regVec_3758 <= _zz_regVec_0;
          end
          if(_zz_1[3759]) begin
            regVec_3759 <= _zz_regVec_0;
          end
          if(_zz_1[3760]) begin
            regVec_3760 <= _zz_regVec_0;
          end
          if(_zz_1[3761]) begin
            regVec_3761 <= _zz_regVec_0;
          end
          if(_zz_1[3762]) begin
            regVec_3762 <= _zz_regVec_0;
          end
          if(_zz_1[3763]) begin
            regVec_3763 <= _zz_regVec_0;
          end
          if(_zz_1[3764]) begin
            regVec_3764 <= _zz_regVec_0;
          end
          if(_zz_1[3765]) begin
            regVec_3765 <= _zz_regVec_0;
          end
          if(_zz_1[3766]) begin
            regVec_3766 <= _zz_regVec_0;
          end
          if(_zz_1[3767]) begin
            regVec_3767 <= _zz_regVec_0;
          end
          if(_zz_1[3768]) begin
            regVec_3768 <= _zz_regVec_0;
          end
          if(_zz_1[3769]) begin
            regVec_3769 <= _zz_regVec_0;
          end
          if(_zz_1[3770]) begin
            regVec_3770 <= _zz_regVec_0;
          end
          if(_zz_1[3771]) begin
            regVec_3771 <= _zz_regVec_0;
          end
          if(_zz_1[3772]) begin
            regVec_3772 <= _zz_regVec_0;
          end
          if(_zz_1[3773]) begin
            regVec_3773 <= _zz_regVec_0;
          end
          if(_zz_1[3774]) begin
            regVec_3774 <= _zz_regVec_0;
          end
          if(_zz_1[3775]) begin
            regVec_3775 <= _zz_regVec_0;
          end
          if(_zz_1[3776]) begin
            regVec_3776 <= _zz_regVec_0;
          end
          if(_zz_1[3777]) begin
            regVec_3777 <= _zz_regVec_0;
          end
          if(_zz_1[3778]) begin
            regVec_3778 <= _zz_regVec_0;
          end
          if(_zz_1[3779]) begin
            regVec_3779 <= _zz_regVec_0;
          end
          if(_zz_1[3780]) begin
            regVec_3780 <= _zz_regVec_0;
          end
          if(_zz_1[3781]) begin
            regVec_3781 <= _zz_regVec_0;
          end
          if(_zz_1[3782]) begin
            regVec_3782 <= _zz_regVec_0;
          end
          if(_zz_1[3783]) begin
            regVec_3783 <= _zz_regVec_0;
          end
          if(_zz_1[3784]) begin
            regVec_3784 <= _zz_regVec_0;
          end
          if(_zz_1[3785]) begin
            regVec_3785 <= _zz_regVec_0;
          end
          if(_zz_1[3786]) begin
            regVec_3786 <= _zz_regVec_0;
          end
          if(_zz_1[3787]) begin
            regVec_3787 <= _zz_regVec_0;
          end
          if(_zz_1[3788]) begin
            regVec_3788 <= _zz_regVec_0;
          end
          if(_zz_1[3789]) begin
            regVec_3789 <= _zz_regVec_0;
          end
          if(_zz_1[3790]) begin
            regVec_3790 <= _zz_regVec_0;
          end
          if(_zz_1[3791]) begin
            regVec_3791 <= _zz_regVec_0;
          end
          if(_zz_1[3792]) begin
            regVec_3792 <= _zz_regVec_0;
          end
          if(_zz_1[3793]) begin
            regVec_3793 <= _zz_regVec_0;
          end
          if(_zz_1[3794]) begin
            regVec_3794 <= _zz_regVec_0;
          end
          if(_zz_1[3795]) begin
            regVec_3795 <= _zz_regVec_0;
          end
          if(_zz_1[3796]) begin
            regVec_3796 <= _zz_regVec_0;
          end
          if(_zz_1[3797]) begin
            regVec_3797 <= _zz_regVec_0;
          end
          if(_zz_1[3798]) begin
            regVec_3798 <= _zz_regVec_0;
          end
          if(_zz_1[3799]) begin
            regVec_3799 <= _zz_regVec_0;
          end
          if(_zz_1[3800]) begin
            regVec_3800 <= _zz_regVec_0;
          end
          if(_zz_1[3801]) begin
            regVec_3801 <= _zz_regVec_0;
          end
          if(_zz_1[3802]) begin
            regVec_3802 <= _zz_regVec_0;
          end
          if(_zz_1[3803]) begin
            regVec_3803 <= _zz_regVec_0;
          end
          if(_zz_1[3804]) begin
            regVec_3804 <= _zz_regVec_0;
          end
          if(_zz_1[3805]) begin
            regVec_3805 <= _zz_regVec_0;
          end
          if(_zz_1[3806]) begin
            regVec_3806 <= _zz_regVec_0;
          end
          if(_zz_1[3807]) begin
            regVec_3807 <= _zz_regVec_0;
          end
          if(_zz_1[3808]) begin
            regVec_3808 <= _zz_regVec_0;
          end
          if(_zz_1[3809]) begin
            regVec_3809 <= _zz_regVec_0;
          end
          if(_zz_1[3810]) begin
            regVec_3810 <= _zz_regVec_0;
          end
          if(_zz_1[3811]) begin
            regVec_3811 <= _zz_regVec_0;
          end
          if(_zz_1[3812]) begin
            regVec_3812 <= _zz_regVec_0;
          end
          if(_zz_1[3813]) begin
            regVec_3813 <= _zz_regVec_0;
          end
          if(_zz_1[3814]) begin
            regVec_3814 <= _zz_regVec_0;
          end
          if(_zz_1[3815]) begin
            regVec_3815 <= _zz_regVec_0;
          end
          if(_zz_1[3816]) begin
            regVec_3816 <= _zz_regVec_0;
          end
          if(_zz_1[3817]) begin
            regVec_3817 <= _zz_regVec_0;
          end
          if(_zz_1[3818]) begin
            regVec_3818 <= _zz_regVec_0;
          end
          if(_zz_1[3819]) begin
            regVec_3819 <= _zz_regVec_0;
          end
          if(_zz_1[3820]) begin
            regVec_3820 <= _zz_regVec_0;
          end
          if(_zz_1[3821]) begin
            regVec_3821 <= _zz_regVec_0;
          end
          if(_zz_1[3822]) begin
            regVec_3822 <= _zz_regVec_0;
          end
          if(_zz_1[3823]) begin
            regVec_3823 <= _zz_regVec_0;
          end
          if(_zz_1[3824]) begin
            regVec_3824 <= _zz_regVec_0;
          end
          if(_zz_1[3825]) begin
            regVec_3825 <= _zz_regVec_0;
          end
          if(_zz_1[3826]) begin
            regVec_3826 <= _zz_regVec_0;
          end
          if(_zz_1[3827]) begin
            regVec_3827 <= _zz_regVec_0;
          end
          if(_zz_1[3828]) begin
            regVec_3828 <= _zz_regVec_0;
          end
          if(_zz_1[3829]) begin
            regVec_3829 <= _zz_regVec_0;
          end
          if(_zz_1[3830]) begin
            regVec_3830 <= _zz_regVec_0;
          end
          if(_zz_1[3831]) begin
            regVec_3831 <= _zz_regVec_0;
          end
          if(_zz_1[3832]) begin
            regVec_3832 <= _zz_regVec_0;
          end
          if(_zz_1[3833]) begin
            regVec_3833 <= _zz_regVec_0;
          end
          if(_zz_1[3834]) begin
            regVec_3834 <= _zz_regVec_0;
          end
          if(_zz_1[3835]) begin
            regVec_3835 <= _zz_regVec_0;
          end
          if(_zz_1[3836]) begin
            regVec_3836 <= _zz_regVec_0;
          end
          if(_zz_1[3837]) begin
            regVec_3837 <= _zz_regVec_0;
          end
          if(_zz_1[3838]) begin
            regVec_3838 <= _zz_regVec_0;
          end
          if(_zz_1[3839]) begin
            regVec_3839 <= _zz_regVec_0;
          end
          if(_zz_1[3840]) begin
            regVec_3840 <= _zz_regVec_0;
          end
          if(_zz_1[3841]) begin
            regVec_3841 <= _zz_regVec_0;
          end
          if(_zz_1[3842]) begin
            regVec_3842 <= _zz_regVec_0;
          end
          if(_zz_1[3843]) begin
            regVec_3843 <= _zz_regVec_0;
          end
          if(_zz_1[3844]) begin
            regVec_3844 <= _zz_regVec_0;
          end
          if(_zz_1[3845]) begin
            regVec_3845 <= _zz_regVec_0;
          end
          if(_zz_1[3846]) begin
            regVec_3846 <= _zz_regVec_0;
          end
          if(_zz_1[3847]) begin
            regVec_3847 <= _zz_regVec_0;
          end
          if(_zz_1[3848]) begin
            regVec_3848 <= _zz_regVec_0;
          end
          if(_zz_1[3849]) begin
            regVec_3849 <= _zz_regVec_0;
          end
          if(_zz_1[3850]) begin
            regVec_3850 <= _zz_regVec_0;
          end
          if(_zz_1[3851]) begin
            regVec_3851 <= _zz_regVec_0;
          end
          if(_zz_1[3852]) begin
            regVec_3852 <= _zz_regVec_0;
          end
          if(_zz_1[3853]) begin
            regVec_3853 <= _zz_regVec_0;
          end
          if(_zz_1[3854]) begin
            regVec_3854 <= _zz_regVec_0;
          end
          if(_zz_1[3855]) begin
            regVec_3855 <= _zz_regVec_0;
          end
          if(_zz_1[3856]) begin
            regVec_3856 <= _zz_regVec_0;
          end
          if(_zz_1[3857]) begin
            regVec_3857 <= _zz_regVec_0;
          end
          if(_zz_1[3858]) begin
            regVec_3858 <= _zz_regVec_0;
          end
          if(_zz_1[3859]) begin
            regVec_3859 <= _zz_regVec_0;
          end
          if(_zz_1[3860]) begin
            regVec_3860 <= _zz_regVec_0;
          end
          if(_zz_1[3861]) begin
            regVec_3861 <= _zz_regVec_0;
          end
          if(_zz_1[3862]) begin
            regVec_3862 <= _zz_regVec_0;
          end
          if(_zz_1[3863]) begin
            regVec_3863 <= _zz_regVec_0;
          end
          if(_zz_1[3864]) begin
            regVec_3864 <= _zz_regVec_0;
          end
          if(_zz_1[3865]) begin
            regVec_3865 <= _zz_regVec_0;
          end
          if(_zz_1[3866]) begin
            regVec_3866 <= _zz_regVec_0;
          end
          if(_zz_1[3867]) begin
            regVec_3867 <= _zz_regVec_0;
          end
          if(_zz_1[3868]) begin
            regVec_3868 <= _zz_regVec_0;
          end
          if(_zz_1[3869]) begin
            regVec_3869 <= _zz_regVec_0;
          end
          if(_zz_1[3870]) begin
            regVec_3870 <= _zz_regVec_0;
          end
          if(_zz_1[3871]) begin
            regVec_3871 <= _zz_regVec_0;
          end
          if(_zz_1[3872]) begin
            regVec_3872 <= _zz_regVec_0;
          end
          if(_zz_1[3873]) begin
            regVec_3873 <= _zz_regVec_0;
          end
          if(_zz_1[3874]) begin
            regVec_3874 <= _zz_regVec_0;
          end
          if(_zz_1[3875]) begin
            regVec_3875 <= _zz_regVec_0;
          end
          if(_zz_1[3876]) begin
            regVec_3876 <= _zz_regVec_0;
          end
          if(_zz_1[3877]) begin
            regVec_3877 <= _zz_regVec_0;
          end
          if(_zz_1[3878]) begin
            regVec_3878 <= _zz_regVec_0;
          end
          if(_zz_1[3879]) begin
            regVec_3879 <= _zz_regVec_0;
          end
          if(_zz_1[3880]) begin
            regVec_3880 <= _zz_regVec_0;
          end
          if(_zz_1[3881]) begin
            regVec_3881 <= _zz_regVec_0;
          end
          if(_zz_1[3882]) begin
            regVec_3882 <= _zz_regVec_0;
          end
          if(_zz_1[3883]) begin
            regVec_3883 <= _zz_regVec_0;
          end
          if(_zz_1[3884]) begin
            regVec_3884 <= _zz_regVec_0;
          end
          if(_zz_1[3885]) begin
            regVec_3885 <= _zz_regVec_0;
          end
          if(_zz_1[3886]) begin
            regVec_3886 <= _zz_regVec_0;
          end
          if(_zz_1[3887]) begin
            regVec_3887 <= _zz_regVec_0;
          end
          if(_zz_1[3888]) begin
            regVec_3888 <= _zz_regVec_0;
          end
          if(_zz_1[3889]) begin
            regVec_3889 <= _zz_regVec_0;
          end
          if(_zz_1[3890]) begin
            regVec_3890 <= _zz_regVec_0;
          end
          if(_zz_1[3891]) begin
            regVec_3891 <= _zz_regVec_0;
          end
          if(_zz_1[3892]) begin
            regVec_3892 <= _zz_regVec_0;
          end
          if(_zz_1[3893]) begin
            regVec_3893 <= _zz_regVec_0;
          end
          if(_zz_1[3894]) begin
            regVec_3894 <= _zz_regVec_0;
          end
          if(_zz_1[3895]) begin
            regVec_3895 <= _zz_regVec_0;
          end
          if(_zz_1[3896]) begin
            regVec_3896 <= _zz_regVec_0;
          end
          if(_zz_1[3897]) begin
            regVec_3897 <= _zz_regVec_0;
          end
          if(_zz_1[3898]) begin
            regVec_3898 <= _zz_regVec_0;
          end
          if(_zz_1[3899]) begin
            regVec_3899 <= _zz_regVec_0;
          end
          if(_zz_1[3900]) begin
            regVec_3900 <= _zz_regVec_0;
          end
          if(_zz_1[3901]) begin
            regVec_3901 <= _zz_regVec_0;
          end
          if(_zz_1[3902]) begin
            regVec_3902 <= _zz_regVec_0;
          end
          if(_zz_1[3903]) begin
            regVec_3903 <= _zz_regVec_0;
          end
          if(_zz_1[3904]) begin
            regVec_3904 <= _zz_regVec_0;
          end
          if(_zz_1[3905]) begin
            regVec_3905 <= _zz_regVec_0;
          end
          if(_zz_1[3906]) begin
            regVec_3906 <= _zz_regVec_0;
          end
          if(_zz_1[3907]) begin
            regVec_3907 <= _zz_regVec_0;
          end
          if(_zz_1[3908]) begin
            regVec_3908 <= _zz_regVec_0;
          end
          if(_zz_1[3909]) begin
            regVec_3909 <= _zz_regVec_0;
          end
          if(_zz_1[3910]) begin
            regVec_3910 <= _zz_regVec_0;
          end
          if(_zz_1[3911]) begin
            regVec_3911 <= _zz_regVec_0;
          end
          if(_zz_1[3912]) begin
            regVec_3912 <= _zz_regVec_0;
          end
          if(_zz_1[3913]) begin
            regVec_3913 <= _zz_regVec_0;
          end
          if(_zz_1[3914]) begin
            regVec_3914 <= _zz_regVec_0;
          end
          if(_zz_1[3915]) begin
            regVec_3915 <= _zz_regVec_0;
          end
          if(_zz_1[3916]) begin
            regVec_3916 <= _zz_regVec_0;
          end
          if(_zz_1[3917]) begin
            regVec_3917 <= _zz_regVec_0;
          end
          if(_zz_1[3918]) begin
            regVec_3918 <= _zz_regVec_0;
          end
          if(_zz_1[3919]) begin
            regVec_3919 <= _zz_regVec_0;
          end
          if(_zz_1[3920]) begin
            regVec_3920 <= _zz_regVec_0;
          end
          if(_zz_1[3921]) begin
            regVec_3921 <= _zz_regVec_0;
          end
          if(_zz_1[3922]) begin
            regVec_3922 <= _zz_regVec_0;
          end
          if(_zz_1[3923]) begin
            regVec_3923 <= _zz_regVec_0;
          end
          if(_zz_1[3924]) begin
            regVec_3924 <= _zz_regVec_0;
          end
          if(_zz_1[3925]) begin
            regVec_3925 <= _zz_regVec_0;
          end
          if(_zz_1[3926]) begin
            regVec_3926 <= _zz_regVec_0;
          end
          if(_zz_1[3927]) begin
            regVec_3927 <= _zz_regVec_0;
          end
          if(_zz_1[3928]) begin
            regVec_3928 <= _zz_regVec_0;
          end
          if(_zz_1[3929]) begin
            regVec_3929 <= _zz_regVec_0;
          end
          if(_zz_1[3930]) begin
            regVec_3930 <= _zz_regVec_0;
          end
          if(_zz_1[3931]) begin
            regVec_3931 <= _zz_regVec_0;
          end
          if(_zz_1[3932]) begin
            regVec_3932 <= _zz_regVec_0;
          end
          if(_zz_1[3933]) begin
            regVec_3933 <= _zz_regVec_0;
          end
          if(_zz_1[3934]) begin
            regVec_3934 <= _zz_regVec_0;
          end
          if(_zz_1[3935]) begin
            regVec_3935 <= _zz_regVec_0;
          end
          if(_zz_1[3936]) begin
            regVec_3936 <= _zz_regVec_0;
          end
          if(_zz_1[3937]) begin
            regVec_3937 <= _zz_regVec_0;
          end
          if(_zz_1[3938]) begin
            regVec_3938 <= _zz_regVec_0;
          end
          if(_zz_1[3939]) begin
            regVec_3939 <= _zz_regVec_0;
          end
          if(_zz_1[3940]) begin
            regVec_3940 <= _zz_regVec_0;
          end
          if(_zz_1[3941]) begin
            regVec_3941 <= _zz_regVec_0;
          end
          if(_zz_1[3942]) begin
            regVec_3942 <= _zz_regVec_0;
          end
          if(_zz_1[3943]) begin
            regVec_3943 <= _zz_regVec_0;
          end
          if(_zz_1[3944]) begin
            regVec_3944 <= _zz_regVec_0;
          end
          if(_zz_1[3945]) begin
            regVec_3945 <= _zz_regVec_0;
          end
          if(_zz_1[3946]) begin
            regVec_3946 <= _zz_regVec_0;
          end
          if(_zz_1[3947]) begin
            regVec_3947 <= _zz_regVec_0;
          end
          if(_zz_1[3948]) begin
            regVec_3948 <= _zz_regVec_0;
          end
          if(_zz_1[3949]) begin
            regVec_3949 <= _zz_regVec_0;
          end
          if(_zz_1[3950]) begin
            regVec_3950 <= _zz_regVec_0;
          end
          if(_zz_1[3951]) begin
            regVec_3951 <= _zz_regVec_0;
          end
          if(_zz_1[3952]) begin
            regVec_3952 <= _zz_regVec_0;
          end
          if(_zz_1[3953]) begin
            regVec_3953 <= _zz_regVec_0;
          end
          if(_zz_1[3954]) begin
            regVec_3954 <= _zz_regVec_0;
          end
          if(_zz_1[3955]) begin
            regVec_3955 <= _zz_regVec_0;
          end
          if(_zz_1[3956]) begin
            regVec_3956 <= _zz_regVec_0;
          end
          if(_zz_1[3957]) begin
            regVec_3957 <= _zz_regVec_0;
          end
          if(_zz_1[3958]) begin
            regVec_3958 <= _zz_regVec_0;
          end
          if(_zz_1[3959]) begin
            regVec_3959 <= _zz_regVec_0;
          end
          if(_zz_1[3960]) begin
            regVec_3960 <= _zz_regVec_0;
          end
          if(_zz_1[3961]) begin
            regVec_3961 <= _zz_regVec_0;
          end
          if(_zz_1[3962]) begin
            regVec_3962 <= _zz_regVec_0;
          end
          if(_zz_1[3963]) begin
            regVec_3963 <= _zz_regVec_0;
          end
          if(_zz_1[3964]) begin
            regVec_3964 <= _zz_regVec_0;
          end
          if(_zz_1[3965]) begin
            regVec_3965 <= _zz_regVec_0;
          end
          if(_zz_1[3966]) begin
            regVec_3966 <= _zz_regVec_0;
          end
          if(_zz_1[3967]) begin
            regVec_3967 <= _zz_regVec_0;
          end
          if(_zz_1[3968]) begin
            regVec_3968 <= _zz_regVec_0;
          end
          if(_zz_1[3969]) begin
            regVec_3969 <= _zz_regVec_0;
          end
          if(_zz_1[3970]) begin
            regVec_3970 <= _zz_regVec_0;
          end
          if(_zz_1[3971]) begin
            regVec_3971 <= _zz_regVec_0;
          end
          if(_zz_1[3972]) begin
            regVec_3972 <= _zz_regVec_0;
          end
          if(_zz_1[3973]) begin
            regVec_3973 <= _zz_regVec_0;
          end
          if(_zz_1[3974]) begin
            regVec_3974 <= _zz_regVec_0;
          end
          if(_zz_1[3975]) begin
            regVec_3975 <= _zz_regVec_0;
          end
          if(_zz_1[3976]) begin
            regVec_3976 <= _zz_regVec_0;
          end
          if(_zz_1[3977]) begin
            regVec_3977 <= _zz_regVec_0;
          end
          if(_zz_1[3978]) begin
            regVec_3978 <= _zz_regVec_0;
          end
          if(_zz_1[3979]) begin
            regVec_3979 <= _zz_regVec_0;
          end
          if(_zz_1[3980]) begin
            regVec_3980 <= _zz_regVec_0;
          end
          if(_zz_1[3981]) begin
            regVec_3981 <= _zz_regVec_0;
          end
          if(_zz_1[3982]) begin
            regVec_3982 <= _zz_regVec_0;
          end
          if(_zz_1[3983]) begin
            regVec_3983 <= _zz_regVec_0;
          end
          if(_zz_1[3984]) begin
            regVec_3984 <= _zz_regVec_0;
          end
          if(_zz_1[3985]) begin
            regVec_3985 <= _zz_regVec_0;
          end
          if(_zz_1[3986]) begin
            regVec_3986 <= _zz_regVec_0;
          end
          if(_zz_1[3987]) begin
            regVec_3987 <= _zz_regVec_0;
          end
          if(_zz_1[3988]) begin
            regVec_3988 <= _zz_regVec_0;
          end
          if(_zz_1[3989]) begin
            regVec_3989 <= _zz_regVec_0;
          end
          if(_zz_1[3990]) begin
            regVec_3990 <= _zz_regVec_0;
          end
          if(_zz_1[3991]) begin
            regVec_3991 <= _zz_regVec_0;
          end
          if(_zz_1[3992]) begin
            regVec_3992 <= _zz_regVec_0;
          end
          if(_zz_1[3993]) begin
            regVec_3993 <= _zz_regVec_0;
          end
          if(_zz_1[3994]) begin
            regVec_3994 <= _zz_regVec_0;
          end
          if(_zz_1[3995]) begin
            regVec_3995 <= _zz_regVec_0;
          end
          if(_zz_1[3996]) begin
            regVec_3996 <= _zz_regVec_0;
          end
          if(_zz_1[3997]) begin
            regVec_3997 <= _zz_regVec_0;
          end
          if(_zz_1[3998]) begin
            regVec_3998 <= _zz_regVec_0;
          end
          if(_zz_1[3999]) begin
            regVec_3999 <= _zz_regVec_0;
          end
          if(_zz_1[4000]) begin
            regVec_4000 <= _zz_regVec_0;
          end
          if(_zz_1[4001]) begin
            regVec_4001 <= _zz_regVec_0;
          end
          if(_zz_1[4002]) begin
            regVec_4002 <= _zz_regVec_0;
          end
          if(_zz_1[4003]) begin
            regVec_4003 <= _zz_regVec_0;
          end
          if(_zz_1[4004]) begin
            regVec_4004 <= _zz_regVec_0;
          end
          if(_zz_1[4005]) begin
            regVec_4005 <= _zz_regVec_0;
          end
          if(_zz_1[4006]) begin
            regVec_4006 <= _zz_regVec_0;
          end
          if(_zz_1[4007]) begin
            regVec_4007 <= _zz_regVec_0;
          end
          if(_zz_1[4008]) begin
            regVec_4008 <= _zz_regVec_0;
          end
          if(_zz_1[4009]) begin
            regVec_4009 <= _zz_regVec_0;
          end
          if(_zz_1[4010]) begin
            regVec_4010 <= _zz_regVec_0;
          end
          if(_zz_1[4011]) begin
            regVec_4011 <= _zz_regVec_0;
          end
          if(_zz_1[4012]) begin
            regVec_4012 <= _zz_regVec_0;
          end
          if(_zz_1[4013]) begin
            regVec_4013 <= _zz_regVec_0;
          end
          if(_zz_1[4014]) begin
            regVec_4014 <= _zz_regVec_0;
          end
          if(_zz_1[4015]) begin
            regVec_4015 <= _zz_regVec_0;
          end
          if(_zz_1[4016]) begin
            regVec_4016 <= _zz_regVec_0;
          end
          if(_zz_1[4017]) begin
            regVec_4017 <= _zz_regVec_0;
          end
          if(_zz_1[4018]) begin
            regVec_4018 <= _zz_regVec_0;
          end
          if(_zz_1[4019]) begin
            regVec_4019 <= _zz_regVec_0;
          end
          if(_zz_1[4020]) begin
            regVec_4020 <= _zz_regVec_0;
          end
          if(_zz_1[4021]) begin
            regVec_4021 <= _zz_regVec_0;
          end
          if(_zz_1[4022]) begin
            regVec_4022 <= _zz_regVec_0;
          end
          if(_zz_1[4023]) begin
            regVec_4023 <= _zz_regVec_0;
          end
          if(_zz_1[4024]) begin
            regVec_4024 <= _zz_regVec_0;
          end
          if(_zz_1[4025]) begin
            regVec_4025 <= _zz_regVec_0;
          end
          if(_zz_1[4026]) begin
            regVec_4026 <= _zz_regVec_0;
          end
          if(_zz_1[4027]) begin
            regVec_4027 <= _zz_regVec_0;
          end
          if(_zz_1[4028]) begin
            regVec_4028 <= _zz_regVec_0;
          end
          if(_zz_1[4029]) begin
            regVec_4029 <= _zz_regVec_0;
          end
          if(_zz_1[4030]) begin
            regVec_4030 <= _zz_regVec_0;
          end
          if(_zz_1[4031]) begin
            regVec_4031 <= _zz_regVec_0;
          end
          if(_zz_1[4032]) begin
            regVec_4032 <= _zz_regVec_0;
          end
          if(_zz_1[4033]) begin
            regVec_4033 <= _zz_regVec_0;
          end
          if(_zz_1[4034]) begin
            regVec_4034 <= _zz_regVec_0;
          end
          if(_zz_1[4035]) begin
            regVec_4035 <= _zz_regVec_0;
          end
          if(_zz_1[4036]) begin
            regVec_4036 <= _zz_regVec_0;
          end
          if(_zz_1[4037]) begin
            regVec_4037 <= _zz_regVec_0;
          end
          if(_zz_1[4038]) begin
            regVec_4038 <= _zz_regVec_0;
          end
          if(_zz_1[4039]) begin
            regVec_4039 <= _zz_regVec_0;
          end
          if(_zz_1[4040]) begin
            regVec_4040 <= _zz_regVec_0;
          end
          if(_zz_1[4041]) begin
            regVec_4041 <= _zz_regVec_0;
          end
          if(_zz_1[4042]) begin
            regVec_4042 <= _zz_regVec_0;
          end
          if(_zz_1[4043]) begin
            regVec_4043 <= _zz_regVec_0;
          end
          if(_zz_1[4044]) begin
            regVec_4044 <= _zz_regVec_0;
          end
          if(_zz_1[4045]) begin
            regVec_4045 <= _zz_regVec_0;
          end
          if(_zz_1[4046]) begin
            regVec_4046 <= _zz_regVec_0;
          end
          if(_zz_1[4047]) begin
            regVec_4047 <= _zz_regVec_0;
          end
          if(_zz_1[4048]) begin
            regVec_4048 <= _zz_regVec_0;
          end
          if(_zz_1[4049]) begin
            regVec_4049 <= _zz_regVec_0;
          end
          if(_zz_1[4050]) begin
            regVec_4050 <= _zz_regVec_0;
          end
          if(_zz_1[4051]) begin
            regVec_4051 <= _zz_regVec_0;
          end
          if(_zz_1[4052]) begin
            regVec_4052 <= _zz_regVec_0;
          end
          if(_zz_1[4053]) begin
            regVec_4053 <= _zz_regVec_0;
          end
          if(_zz_1[4054]) begin
            regVec_4054 <= _zz_regVec_0;
          end
          if(_zz_1[4055]) begin
            regVec_4055 <= _zz_regVec_0;
          end
          if(_zz_1[4056]) begin
            regVec_4056 <= _zz_regVec_0;
          end
          if(_zz_1[4057]) begin
            regVec_4057 <= _zz_regVec_0;
          end
          if(_zz_1[4058]) begin
            regVec_4058 <= _zz_regVec_0;
          end
          if(_zz_1[4059]) begin
            regVec_4059 <= _zz_regVec_0;
          end
          if(_zz_1[4060]) begin
            regVec_4060 <= _zz_regVec_0;
          end
          if(_zz_1[4061]) begin
            regVec_4061 <= _zz_regVec_0;
          end
          if(_zz_1[4062]) begin
            regVec_4062 <= _zz_regVec_0;
          end
          if(_zz_1[4063]) begin
            regVec_4063 <= _zz_regVec_0;
          end
          if(_zz_1[4064]) begin
            regVec_4064 <= _zz_regVec_0;
          end
          if(_zz_1[4065]) begin
            regVec_4065 <= _zz_regVec_0;
          end
          if(_zz_1[4066]) begin
            regVec_4066 <= _zz_regVec_0;
          end
          if(_zz_1[4067]) begin
            regVec_4067 <= _zz_regVec_0;
          end
          if(_zz_1[4068]) begin
            regVec_4068 <= _zz_regVec_0;
          end
          if(_zz_1[4069]) begin
            regVec_4069 <= _zz_regVec_0;
          end
          if(_zz_1[4070]) begin
            regVec_4070 <= _zz_regVec_0;
          end
          if(_zz_1[4071]) begin
            regVec_4071 <= _zz_regVec_0;
          end
          if(_zz_1[4072]) begin
            regVec_4072 <= _zz_regVec_0;
          end
          if(_zz_1[4073]) begin
            regVec_4073 <= _zz_regVec_0;
          end
          if(_zz_1[4074]) begin
            regVec_4074 <= _zz_regVec_0;
          end
          if(_zz_1[4075]) begin
            regVec_4075 <= _zz_regVec_0;
          end
          if(_zz_1[4076]) begin
            regVec_4076 <= _zz_regVec_0;
          end
          if(_zz_1[4077]) begin
            regVec_4077 <= _zz_regVec_0;
          end
          if(_zz_1[4078]) begin
            regVec_4078 <= _zz_regVec_0;
          end
          if(_zz_1[4079]) begin
            regVec_4079 <= _zz_regVec_0;
          end
          if(_zz_1[4080]) begin
            regVec_4080 <= _zz_regVec_0;
          end
          if(_zz_1[4081]) begin
            regVec_4081 <= _zz_regVec_0;
          end
          if(_zz_1[4082]) begin
            regVec_4082 <= _zz_regVec_0;
          end
          if(_zz_1[4083]) begin
            regVec_4083 <= _zz_regVec_0;
          end
          if(_zz_1[4084]) begin
            regVec_4084 <= _zz_regVec_0;
          end
          if(_zz_1[4085]) begin
            regVec_4085 <= _zz_regVec_0;
          end
          if(_zz_1[4086]) begin
            regVec_4086 <= _zz_regVec_0;
          end
          if(_zz_1[4087]) begin
            regVec_4087 <= _zz_regVec_0;
          end
          if(_zz_1[4088]) begin
            regVec_4088 <= _zz_regVec_0;
          end
          if(_zz_1[4089]) begin
            regVec_4089 <= _zz_regVec_0;
          end
          if(_zz_1[4090]) begin
            regVec_4090 <= _zz_regVec_0;
          end
          if(_zz_1[4091]) begin
            regVec_4091 <= _zz_regVec_0;
          end
          if(_zz_1[4092]) begin
            regVec_4092 <= _zz_regVec_0;
          end
          if(_zz_1[4093]) begin
            regVec_4093 <= _zz_regVec_0;
          end
          if(_zz_1[4094]) begin
            regVec_4094 <= _zz_regVec_0;
          end
          if(_zz_1[4095]) begin
            regVec_4095 <= _zz_regVec_0;
          end
        end else begin
          if(_zz_2[0]) begin
            regVec_0 <= _zz_regVec_0_1;
          end
          if(_zz_2[1]) begin
            regVec_1 <= _zz_regVec_0_1;
          end
          if(_zz_2[2]) begin
            regVec_2 <= _zz_regVec_0_1;
          end
          if(_zz_2[3]) begin
            regVec_3 <= _zz_regVec_0_1;
          end
          if(_zz_2[4]) begin
            regVec_4 <= _zz_regVec_0_1;
          end
          if(_zz_2[5]) begin
            regVec_5 <= _zz_regVec_0_1;
          end
          if(_zz_2[6]) begin
            regVec_6 <= _zz_regVec_0_1;
          end
          if(_zz_2[7]) begin
            regVec_7 <= _zz_regVec_0_1;
          end
          if(_zz_2[8]) begin
            regVec_8 <= _zz_regVec_0_1;
          end
          if(_zz_2[9]) begin
            regVec_9 <= _zz_regVec_0_1;
          end
          if(_zz_2[10]) begin
            regVec_10 <= _zz_regVec_0_1;
          end
          if(_zz_2[11]) begin
            regVec_11 <= _zz_regVec_0_1;
          end
          if(_zz_2[12]) begin
            regVec_12 <= _zz_regVec_0_1;
          end
          if(_zz_2[13]) begin
            regVec_13 <= _zz_regVec_0_1;
          end
          if(_zz_2[14]) begin
            regVec_14 <= _zz_regVec_0_1;
          end
          if(_zz_2[15]) begin
            regVec_15 <= _zz_regVec_0_1;
          end
          if(_zz_2[16]) begin
            regVec_16 <= _zz_regVec_0_1;
          end
          if(_zz_2[17]) begin
            regVec_17 <= _zz_regVec_0_1;
          end
          if(_zz_2[18]) begin
            regVec_18 <= _zz_regVec_0_1;
          end
          if(_zz_2[19]) begin
            regVec_19 <= _zz_regVec_0_1;
          end
          if(_zz_2[20]) begin
            regVec_20 <= _zz_regVec_0_1;
          end
          if(_zz_2[21]) begin
            regVec_21 <= _zz_regVec_0_1;
          end
          if(_zz_2[22]) begin
            regVec_22 <= _zz_regVec_0_1;
          end
          if(_zz_2[23]) begin
            regVec_23 <= _zz_regVec_0_1;
          end
          if(_zz_2[24]) begin
            regVec_24 <= _zz_regVec_0_1;
          end
          if(_zz_2[25]) begin
            regVec_25 <= _zz_regVec_0_1;
          end
          if(_zz_2[26]) begin
            regVec_26 <= _zz_regVec_0_1;
          end
          if(_zz_2[27]) begin
            regVec_27 <= _zz_regVec_0_1;
          end
          if(_zz_2[28]) begin
            regVec_28 <= _zz_regVec_0_1;
          end
          if(_zz_2[29]) begin
            regVec_29 <= _zz_regVec_0_1;
          end
          if(_zz_2[30]) begin
            regVec_30 <= _zz_regVec_0_1;
          end
          if(_zz_2[31]) begin
            regVec_31 <= _zz_regVec_0_1;
          end
          if(_zz_2[32]) begin
            regVec_32 <= _zz_regVec_0_1;
          end
          if(_zz_2[33]) begin
            regVec_33 <= _zz_regVec_0_1;
          end
          if(_zz_2[34]) begin
            regVec_34 <= _zz_regVec_0_1;
          end
          if(_zz_2[35]) begin
            regVec_35 <= _zz_regVec_0_1;
          end
          if(_zz_2[36]) begin
            regVec_36 <= _zz_regVec_0_1;
          end
          if(_zz_2[37]) begin
            regVec_37 <= _zz_regVec_0_1;
          end
          if(_zz_2[38]) begin
            regVec_38 <= _zz_regVec_0_1;
          end
          if(_zz_2[39]) begin
            regVec_39 <= _zz_regVec_0_1;
          end
          if(_zz_2[40]) begin
            regVec_40 <= _zz_regVec_0_1;
          end
          if(_zz_2[41]) begin
            regVec_41 <= _zz_regVec_0_1;
          end
          if(_zz_2[42]) begin
            regVec_42 <= _zz_regVec_0_1;
          end
          if(_zz_2[43]) begin
            regVec_43 <= _zz_regVec_0_1;
          end
          if(_zz_2[44]) begin
            regVec_44 <= _zz_regVec_0_1;
          end
          if(_zz_2[45]) begin
            regVec_45 <= _zz_regVec_0_1;
          end
          if(_zz_2[46]) begin
            regVec_46 <= _zz_regVec_0_1;
          end
          if(_zz_2[47]) begin
            regVec_47 <= _zz_regVec_0_1;
          end
          if(_zz_2[48]) begin
            regVec_48 <= _zz_regVec_0_1;
          end
          if(_zz_2[49]) begin
            regVec_49 <= _zz_regVec_0_1;
          end
          if(_zz_2[50]) begin
            regVec_50 <= _zz_regVec_0_1;
          end
          if(_zz_2[51]) begin
            regVec_51 <= _zz_regVec_0_1;
          end
          if(_zz_2[52]) begin
            regVec_52 <= _zz_regVec_0_1;
          end
          if(_zz_2[53]) begin
            regVec_53 <= _zz_regVec_0_1;
          end
          if(_zz_2[54]) begin
            regVec_54 <= _zz_regVec_0_1;
          end
          if(_zz_2[55]) begin
            regVec_55 <= _zz_regVec_0_1;
          end
          if(_zz_2[56]) begin
            regVec_56 <= _zz_regVec_0_1;
          end
          if(_zz_2[57]) begin
            regVec_57 <= _zz_regVec_0_1;
          end
          if(_zz_2[58]) begin
            regVec_58 <= _zz_regVec_0_1;
          end
          if(_zz_2[59]) begin
            regVec_59 <= _zz_regVec_0_1;
          end
          if(_zz_2[60]) begin
            regVec_60 <= _zz_regVec_0_1;
          end
          if(_zz_2[61]) begin
            regVec_61 <= _zz_regVec_0_1;
          end
          if(_zz_2[62]) begin
            regVec_62 <= _zz_regVec_0_1;
          end
          if(_zz_2[63]) begin
            regVec_63 <= _zz_regVec_0_1;
          end
          if(_zz_2[64]) begin
            regVec_64 <= _zz_regVec_0_1;
          end
          if(_zz_2[65]) begin
            regVec_65 <= _zz_regVec_0_1;
          end
          if(_zz_2[66]) begin
            regVec_66 <= _zz_regVec_0_1;
          end
          if(_zz_2[67]) begin
            regVec_67 <= _zz_regVec_0_1;
          end
          if(_zz_2[68]) begin
            regVec_68 <= _zz_regVec_0_1;
          end
          if(_zz_2[69]) begin
            regVec_69 <= _zz_regVec_0_1;
          end
          if(_zz_2[70]) begin
            regVec_70 <= _zz_regVec_0_1;
          end
          if(_zz_2[71]) begin
            regVec_71 <= _zz_regVec_0_1;
          end
          if(_zz_2[72]) begin
            regVec_72 <= _zz_regVec_0_1;
          end
          if(_zz_2[73]) begin
            regVec_73 <= _zz_regVec_0_1;
          end
          if(_zz_2[74]) begin
            regVec_74 <= _zz_regVec_0_1;
          end
          if(_zz_2[75]) begin
            regVec_75 <= _zz_regVec_0_1;
          end
          if(_zz_2[76]) begin
            regVec_76 <= _zz_regVec_0_1;
          end
          if(_zz_2[77]) begin
            regVec_77 <= _zz_regVec_0_1;
          end
          if(_zz_2[78]) begin
            regVec_78 <= _zz_regVec_0_1;
          end
          if(_zz_2[79]) begin
            regVec_79 <= _zz_regVec_0_1;
          end
          if(_zz_2[80]) begin
            regVec_80 <= _zz_regVec_0_1;
          end
          if(_zz_2[81]) begin
            regVec_81 <= _zz_regVec_0_1;
          end
          if(_zz_2[82]) begin
            regVec_82 <= _zz_regVec_0_1;
          end
          if(_zz_2[83]) begin
            regVec_83 <= _zz_regVec_0_1;
          end
          if(_zz_2[84]) begin
            regVec_84 <= _zz_regVec_0_1;
          end
          if(_zz_2[85]) begin
            regVec_85 <= _zz_regVec_0_1;
          end
          if(_zz_2[86]) begin
            regVec_86 <= _zz_regVec_0_1;
          end
          if(_zz_2[87]) begin
            regVec_87 <= _zz_regVec_0_1;
          end
          if(_zz_2[88]) begin
            regVec_88 <= _zz_regVec_0_1;
          end
          if(_zz_2[89]) begin
            regVec_89 <= _zz_regVec_0_1;
          end
          if(_zz_2[90]) begin
            regVec_90 <= _zz_regVec_0_1;
          end
          if(_zz_2[91]) begin
            regVec_91 <= _zz_regVec_0_1;
          end
          if(_zz_2[92]) begin
            regVec_92 <= _zz_regVec_0_1;
          end
          if(_zz_2[93]) begin
            regVec_93 <= _zz_regVec_0_1;
          end
          if(_zz_2[94]) begin
            regVec_94 <= _zz_regVec_0_1;
          end
          if(_zz_2[95]) begin
            regVec_95 <= _zz_regVec_0_1;
          end
          if(_zz_2[96]) begin
            regVec_96 <= _zz_regVec_0_1;
          end
          if(_zz_2[97]) begin
            regVec_97 <= _zz_regVec_0_1;
          end
          if(_zz_2[98]) begin
            regVec_98 <= _zz_regVec_0_1;
          end
          if(_zz_2[99]) begin
            regVec_99 <= _zz_regVec_0_1;
          end
          if(_zz_2[100]) begin
            regVec_100 <= _zz_regVec_0_1;
          end
          if(_zz_2[101]) begin
            regVec_101 <= _zz_regVec_0_1;
          end
          if(_zz_2[102]) begin
            regVec_102 <= _zz_regVec_0_1;
          end
          if(_zz_2[103]) begin
            regVec_103 <= _zz_regVec_0_1;
          end
          if(_zz_2[104]) begin
            regVec_104 <= _zz_regVec_0_1;
          end
          if(_zz_2[105]) begin
            regVec_105 <= _zz_regVec_0_1;
          end
          if(_zz_2[106]) begin
            regVec_106 <= _zz_regVec_0_1;
          end
          if(_zz_2[107]) begin
            regVec_107 <= _zz_regVec_0_1;
          end
          if(_zz_2[108]) begin
            regVec_108 <= _zz_regVec_0_1;
          end
          if(_zz_2[109]) begin
            regVec_109 <= _zz_regVec_0_1;
          end
          if(_zz_2[110]) begin
            regVec_110 <= _zz_regVec_0_1;
          end
          if(_zz_2[111]) begin
            regVec_111 <= _zz_regVec_0_1;
          end
          if(_zz_2[112]) begin
            regVec_112 <= _zz_regVec_0_1;
          end
          if(_zz_2[113]) begin
            regVec_113 <= _zz_regVec_0_1;
          end
          if(_zz_2[114]) begin
            regVec_114 <= _zz_regVec_0_1;
          end
          if(_zz_2[115]) begin
            regVec_115 <= _zz_regVec_0_1;
          end
          if(_zz_2[116]) begin
            regVec_116 <= _zz_regVec_0_1;
          end
          if(_zz_2[117]) begin
            regVec_117 <= _zz_regVec_0_1;
          end
          if(_zz_2[118]) begin
            regVec_118 <= _zz_regVec_0_1;
          end
          if(_zz_2[119]) begin
            regVec_119 <= _zz_regVec_0_1;
          end
          if(_zz_2[120]) begin
            regVec_120 <= _zz_regVec_0_1;
          end
          if(_zz_2[121]) begin
            regVec_121 <= _zz_regVec_0_1;
          end
          if(_zz_2[122]) begin
            regVec_122 <= _zz_regVec_0_1;
          end
          if(_zz_2[123]) begin
            regVec_123 <= _zz_regVec_0_1;
          end
          if(_zz_2[124]) begin
            regVec_124 <= _zz_regVec_0_1;
          end
          if(_zz_2[125]) begin
            regVec_125 <= _zz_regVec_0_1;
          end
          if(_zz_2[126]) begin
            regVec_126 <= _zz_regVec_0_1;
          end
          if(_zz_2[127]) begin
            regVec_127 <= _zz_regVec_0_1;
          end
          if(_zz_2[128]) begin
            regVec_128 <= _zz_regVec_0_1;
          end
          if(_zz_2[129]) begin
            regVec_129 <= _zz_regVec_0_1;
          end
          if(_zz_2[130]) begin
            regVec_130 <= _zz_regVec_0_1;
          end
          if(_zz_2[131]) begin
            regVec_131 <= _zz_regVec_0_1;
          end
          if(_zz_2[132]) begin
            regVec_132 <= _zz_regVec_0_1;
          end
          if(_zz_2[133]) begin
            regVec_133 <= _zz_regVec_0_1;
          end
          if(_zz_2[134]) begin
            regVec_134 <= _zz_regVec_0_1;
          end
          if(_zz_2[135]) begin
            regVec_135 <= _zz_regVec_0_1;
          end
          if(_zz_2[136]) begin
            regVec_136 <= _zz_regVec_0_1;
          end
          if(_zz_2[137]) begin
            regVec_137 <= _zz_regVec_0_1;
          end
          if(_zz_2[138]) begin
            regVec_138 <= _zz_regVec_0_1;
          end
          if(_zz_2[139]) begin
            regVec_139 <= _zz_regVec_0_1;
          end
          if(_zz_2[140]) begin
            regVec_140 <= _zz_regVec_0_1;
          end
          if(_zz_2[141]) begin
            regVec_141 <= _zz_regVec_0_1;
          end
          if(_zz_2[142]) begin
            regVec_142 <= _zz_regVec_0_1;
          end
          if(_zz_2[143]) begin
            regVec_143 <= _zz_regVec_0_1;
          end
          if(_zz_2[144]) begin
            regVec_144 <= _zz_regVec_0_1;
          end
          if(_zz_2[145]) begin
            regVec_145 <= _zz_regVec_0_1;
          end
          if(_zz_2[146]) begin
            regVec_146 <= _zz_regVec_0_1;
          end
          if(_zz_2[147]) begin
            regVec_147 <= _zz_regVec_0_1;
          end
          if(_zz_2[148]) begin
            regVec_148 <= _zz_regVec_0_1;
          end
          if(_zz_2[149]) begin
            regVec_149 <= _zz_regVec_0_1;
          end
          if(_zz_2[150]) begin
            regVec_150 <= _zz_regVec_0_1;
          end
          if(_zz_2[151]) begin
            regVec_151 <= _zz_regVec_0_1;
          end
          if(_zz_2[152]) begin
            regVec_152 <= _zz_regVec_0_1;
          end
          if(_zz_2[153]) begin
            regVec_153 <= _zz_regVec_0_1;
          end
          if(_zz_2[154]) begin
            regVec_154 <= _zz_regVec_0_1;
          end
          if(_zz_2[155]) begin
            regVec_155 <= _zz_regVec_0_1;
          end
          if(_zz_2[156]) begin
            regVec_156 <= _zz_regVec_0_1;
          end
          if(_zz_2[157]) begin
            regVec_157 <= _zz_regVec_0_1;
          end
          if(_zz_2[158]) begin
            regVec_158 <= _zz_regVec_0_1;
          end
          if(_zz_2[159]) begin
            regVec_159 <= _zz_regVec_0_1;
          end
          if(_zz_2[160]) begin
            regVec_160 <= _zz_regVec_0_1;
          end
          if(_zz_2[161]) begin
            regVec_161 <= _zz_regVec_0_1;
          end
          if(_zz_2[162]) begin
            regVec_162 <= _zz_regVec_0_1;
          end
          if(_zz_2[163]) begin
            regVec_163 <= _zz_regVec_0_1;
          end
          if(_zz_2[164]) begin
            regVec_164 <= _zz_regVec_0_1;
          end
          if(_zz_2[165]) begin
            regVec_165 <= _zz_regVec_0_1;
          end
          if(_zz_2[166]) begin
            regVec_166 <= _zz_regVec_0_1;
          end
          if(_zz_2[167]) begin
            regVec_167 <= _zz_regVec_0_1;
          end
          if(_zz_2[168]) begin
            regVec_168 <= _zz_regVec_0_1;
          end
          if(_zz_2[169]) begin
            regVec_169 <= _zz_regVec_0_1;
          end
          if(_zz_2[170]) begin
            regVec_170 <= _zz_regVec_0_1;
          end
          if(_zz_2[171]) begin
            regVec_171 <= _zz_regVec_0_1;
          end
          if(_zz_2[172]) begin
            regVec_172 <= _zz_regVec_0_1;
          end
          if(_zz_2[173]) begin
            regVec_173 <= _zz_regVec_0_1;
          end
          if(_zz_2[174]) begin
            regVec_174 <= _zz_regVec_0_1;
          end
          if(_zz_2[175]) begin
            regVec_175 <= _zz_regVec_0_1;
          end
          if(_zz_2[176]) begin
            regVec_176 <= _zz_regVec_0_1;
          end
          if(_zz_2[177]) begin
            regVec_177 <= _zz_regVec_0_1;
          end
          if(_zz_2[178]) begin
            regVec_178 <= _zz_regVec_0_1;
          end
          if(_zz_2[179]) begin
            regVec_179 <= _zz_regVec_0_1;
          end
          if(_zz_2[180]) begin
            regVec_180 <= _zz_regVec_0_1;
          end
          if(_zz_2[181]) begin
            regVec_181 <= _zz_regVec_0_1;
          end
          if(_zz_2[182]) begin
            regVec_182 <= _zz_regVec_0_1;
          end
          if(_zz_2[183]) begin
            regVec_183 <= _zz_regVec_0_1;
          end
          if(_zz_2[184]) begin
            regVec_184 <= _zz_regVec_0_1;
          end
          if(_zz_2[185]) begin
            regVec_185 <= _zz_regVec_0_1;
          end
          if(_zz_2[186]) begin
            regVec_186 <= _zz_regVec_0_1;
          end
          if(_zz_2[187]) begin
            regVec_187 <= _zz_regVec_0_1;
          end
          if(_zz_2[188]) begin
            regVec_188 <= _zz_regVec_0_1;
          end
          if(_zz_2[189]) begin
            regVec_189 <= _zz_regVec_0_1;
          end
          if(_zz_2[190]) begin
            regVec_190 <= _zz_regVec_0_1;
          end
          if(_zz_2[191]) begin
            regVec_191 <= _zz_regVec_0_1;
          end
          if(_zz_2[192]) begin
            regVec_192 <= _zz_regVec_0_1;
          end
          if(_zz_2[193]) begin
            regVec_193 <= _zz_regVec_0_1;
          end
          if(_zz_2[194]) begin
            regVec_194 <= _zz_regVec_0_1;
          end
          if(_zz_2[195]) begin
            regVec_195 <= _zz_regVec_0_1;
          end
          if(_zz_2[196]) begin
            regVec_196 <= _zz_regVec_0_1;
          end
          if(_zz_2[197]) begin
            regVec_197 <= _zz_regVec_0_1;
          end
          if(_zz_2[198]) begin
            regVec_198 <= _zz_regVec_0_1;
          end
          if(_zz_2[199]) begin
            regVec_199 <= _zz_regVec_0_1;
          end
          if(_zz_2[200]) begin
            regVec_200 <= _zz_regVec_0_1;
          end
          if(_zz_2[201]) begin
            regVec_201 <= _zz_regVec_0_1;
          end
          if(_zz_2[202]) begin
            regVec_202 <= _zz_regVec_0_1;
          end
          if(_zz_2[203]) begin
            regVec_203 <= _zz_regVec_0_1;
          end
          if(_zz_2[204]) begin
            regVec_204 <= _zz_regVec_0_1;
          end
          if(_zz_2[205]) begin
            regVec_205 <= _zz_regVec_0_1;
          end
          if(_zz_2[206]) begin
            regVec_206 <= _zz_regVec_0_1;
          end
          if(_zz_2[207]) begin
            regVec_207 <= _zz_regVec_0_1;
          end
          if(_zz_2[208]) begin
            regVec_208 <= _zz_regVec_0_1;
          end
          if(_zz_2[209]) begin
            regVec_209 <= _zz_regVec_0_1;
          end
          if(_zz_2[210]) begin
            regVec_210 <= _zz_regVec_0_1;
          end
          if(_zz_2[211]) begin
            regVec_211 <= _zz_regVec_0_1;
          end
          if(_zz_2[212]) begin
            regVec_212 <= _zz_regVec_0_1;
          end
          if(_zz_2[213]) begin
            regVec_213 <= _zz_regVec_0_1;
          end
          if(_zz_2[214]) begin
            regVec_214 <= _zz_regVec_0_1;
          end
          if(_zz_2[215]) begin
            regVec_215 <= _zz_regVec_0_1;
          end
          if(_zz_2[216]) begin
            regVec_216 <= _zz_regVec_0_1;
          end
          if(_zz_2[217]) begin
            regVec_217 <= _zz_regVec_0_1;
          end
          if(_zz_2[218]) begin
            regVec_218 <= _zz_regVec_0_1;
          end
          if(_zz_2[219]) begin
            regVec_219 <= _zz_regVec_0_1;
          end
          if(_zz_2[220]) begin
            regVec_220 <= _zz_regVec_0_1;
          end
          if(_zz_2[221]) begin
            regVec_221 <= _zz_regVec_0_1;
          end
          if(_zz_2[222]) begin
            regVec_222 <= _zz_regVec_0_1;
          end
          if(_zz_2[223]) begin
            regVec_223 <= _zz_regVec_0_1;
          end
          if(_zz_2[224]) begin
            regVec_224 <= _zz_regVec_0_1;
          end
          if(_zz_2[225]) begin
            regVec_225 <= _zz_regVec_0_1;
          end
          if(_zz_2[226]) begin
            regVec_226 <= _zz_regVec_0_1;
          end
          if(_zz_2[227]) begin
            regVec_227 <= _zz_regVec_0_1;
          end
          if(_zz_2[228]) begin
            regVec_228 <= _zz_regVec_0_1;
          end
          if(_zz_2[229]) begin
            regVec_229 <= _zz_regVec_0_1;
          end
          if(_zz_2[230]) begin
            regVec_230 <= _zz_regVec_0_1;
          end
          if(_zz_2[231]) begin
            regVec_231 <= _zz_regVec_0_1;
          end
          if(_zz_2[232]) begin
            regVec_232 <= _zz_regVec_0_1;
          end
          if(_zz_2[233]) begin
            regVec_233 <= _zz_regVec_0_1;
          end
          if(_zz_2[234]) begin
            regVec_234 <= _zz_regVec_0_1;
          end
          if(_zz_2[235]) begin
            regVec_235 <= _zz_regVec_0_1;
          end
          if(_zz_2[236]) begin
            regVec_236 <= _zz_regVec_0_1;
          end
          if(_zz_2[237]) begin
            regVec_237 <= _zz_regVec_0_1;
          end
          if(_zz_2[238]) begin
            regVec_238 <= _zz_regVec_0_1;
          end
          if(_zz_2[239]) begin
            regVec_239 <= _zz_regVec_0_1;
          end
          if(_zz_2[240]) begin
            regVec_240 <= _zz_regVec_0_1;
          end
          if(_zz_2[241]) begin
            regVec_241 <= _zz_regVec_0_1;
          end
          if(_zz_2[242]) begin
            regVec_242 <= _zz_regVec_0_1;
          end
          if(_zz_2[243]) begin
            regVec_243 <= _zz_regVec_0_1;
          end
          if(_zz_2[244]) begin
            regVec_244 <= _zz_regVec_0_1;
          end
          if(_zz_2[245]) begin
            regVec_245 <= _zz_regVec_0_1;
          end
          if(_zz_2[246]) begin
            regVec_246 <= _zz_regVec_0_1;
          end
          if(_zz_2[247]) begin
            regVec_247 <= _zz_regVec_0_1;
          end
          if(_zz_2[248]) begin
            regVec_248 <= _zz_regVec_0_1;
          end
          if(_zz_2[249]) begin
            regVec_249 <= _zz_regVec_0_1;
          end
          if(_zz_2[250]) begin
            regVec_250 <= _zz_regVec_0_1;
          end
          if(_zz_2[251]) begin
            regVec_251 <= _zz_regVec_0_1;
          end
          if(_zz_2[252]) begin
            regVec_252 <= _zz_regVec_0_1;
          end
          if(_zz_2[253]) begin
            regVec_253 <= _zz_regVec_0_1;
          end
          if(_zz_2[254]) begin
            regVec_254 <= _zz_regVec_0_1;
          end
          if(_zz_2[255]) begin
            regVec_255 <= _zz_regVec_0_1;
          end
          if(_zz_2[256]) begin
            regVec_256 <= _zz_regVec_0_1;
          end
          if(_zz_2[257]) begin
            regVec_257 <= _zz_regVec_0_1;
          end
          if(_zz_2[258]) begin
            regVec_258 <= _zz_regVec_0_1;
          end
          if(_zz_2[259]) begin
            regVec_259 <= _zz_regVec_0_1;
          end
          if(_zz_2[260]) begin
            regVec_260 <= _zz_regVec_0_1;
          end
          if(_zz_2[261]) begin
            regVec_261 <= _zz_regVec_0_1;
          end
          if(_zz_2[262]) begin
            regVec_262 <= _zz_regVec_0_1;
          end
          if(_zz_2[263]) begin
            regVec_263 <= _zz_regVec_0_1;
          end
          if(_zz_2[264]) begin
            regVec_264 <= _zz_regVec_0_1;
          end
          if(_zz_2[265]) begin
            regVec_265 <= _zz_regVec_0_1;
          end
          if(_zz_2[266]) begin
            regVec_266 <= _zz_regVec_0_1;
          end
          if(_zz_2[267]) begin
            regVec_267 <= _zz_regVec_0_1;
          end
          if(_zz_2[268]) begin
            regVec_268 <= _zz_regVec_0_1;
          end
          if(_zz_2[269]) begin
            regVec_269 <= _zz_regVec_0_1;
          end
          if(_zz_2[270]) begin
            regVec_270 <= _zz_regVec_0_1;
          end
          if(_zz_2[271]) begin
            regVec_271 <= _zz_regVec_0_1;
          end
          if(_zz_2[272]) begin
            regVec_272 <= _zz_regVec_0_1;
          end
          if(_zz_2[273]) begin
            regVec_273 <= _zz_regVec_0_1;
          end
          if(_zz_2[274]) begin
            regVec_274 <= _zz_regVec_0_1;
          end
          if(_zz_2[275]) begin
            regVec_275 <= _zz_regVec_0_1;
          end
          if(_zz_2[276]) begin
            regVec_276 <= _zz_regVec_0_1;
          end
          if(_zz_2[277]) begin
            regVec_277 <= _zz_regVec_0_1;
          end
          if(_zz_2[278]) begin
            regVec_278 <= _zz_regVec_0_1;
          end
          if(_zz_2[279]) begin
            regVec_279 <= _zz_regVec_0_1;
          end
          if(_zz_2[280]) begin
            regVec_280 <= _zz_regVec_0_1;
          end
          if(_zz_2[281]) begin
            regVec_281 <= _zz_regVec_0_1;
          end
          if(_zz_2[282]) begin
            regVec_282 <= _zz_regVec_0_1;
          end
          if(_zz_2[283]) begin
            regVec_283 <= _zz_regVec_0_1;
          end
          if(_zz_2[284]) begin
            regVec_284 <= _zz_regVec_0_1;
          end
          if(_zz_2[285]) begin
            regVec_285 <= _zz_regVec_0_1;
          end
          if(_zz_2[286]) begin
            regVec_286 <= _zz_regVec_0_1;
          end
          if(_zz_2[287]) begin
            regVec_287 <= _zz_regVec_0_1;
          end
          if(_zz_2[288]) begin
            regVec_288 <= _zz_regVec_0_1;
          end
          if(_zz_2[289]) begin
            regVec_289 <= _zz_regVec_0_1;
          end
          if(_zz_2[290]) begin
            regVec_290 <= _zz_regVec_0_1;
          end
          if(_zz_2[291]) begin
            regVec_291 <= _zz_regVec_0_1;
          end
          if(_zz_2[292]) begin
            regVec_292 <= _zz_regVec_0_1;
          end
          if(_zz_2[293]) begin
            regVec_293 <= _zz_regVec_0_1;
          end
          if(_zz_2[294]) begin
            regVec_294 <= _zz_regVec_0_1;
          end
          if(_zz_2[295]) begin
            regVec_295 <= _zz_regVec_0_1;
          end
          if(_zz_2[296]) begin
            regVec_296 <= _zz_regVec_0_1;
          end
          if(_zz_2[297]) begin
            regVec_297 <= _zz_regVec_0_1;
          end
          if(_zz_2[298]) begin
            regVec_298 <= _zz_regVec_0_1;
          end
          if(_zz_2[299]) begin
            regVec_299 <= _zz_regVec_0_1;
          end
          if(_zz_2[300]) begin
            regVec_300 <= _zz_regVec_0_1;
          end
          if(_zz_2[301]) begin
            regVec_301 <= _zz_regVec_0_1;
          end
          if(_zz_2[302]) begin
            regVec_302 <= _zz_regVec_0_1;
          end
          if(_zz_2[303]) begin
            regVec_303 <= _zz_regVec_0_1;
          end
          if(_zz_2[304]) begin
            regVec_304 <= _zz_regVec_0_1;
          end
          if(_zz_2[305]) begin
            regVec_305 <= _zz_regVec_0_1;
          end
          if(_zz_2[306]) begin
            regVec_306 <= _zz_regVec_0_1;
          end
          if(_zz_2[307]) begin
            regVec_307 <= _zz_regVec_0_1;
          end
          if(_zz_2[308]) begin
            regVec_308 <= _zz_regVec_0_1;
          end
          if(_zz_2[309]) begin
            regVec_309 <= _zz_regVec_0_1;
          end
          if(_zz_2[310]) begin
            regVec_310 <= _zz_regVec_0_1;
          end
          if(_zz_2[311]) begin
            regVec_311 <= _zz_regVec_0_1;
          end
          if(_zz_2[312]) begin
            regVec_312 <= _zz_regVec_0_1;
          end
          if(_zz_2[313]) begin
            regVec_313 <= _zz_regVec_0_1;
          end
          if(_zz_2[314]) begin
            regVec_314 <= _zz_regVec_0_1;
          end
          if(_zz_2[315]) begin
            regVec_315 <= _zz_regVec_0_1;
          end
          if(_zz_2[316]) begin
            regVec_316 <= _zz_regVec_0_1;
          end
          if(_zz_2[317]) begin
            regVec_317 <= _zz_regVec_0_1;
          end
          if(_zz_2[318]) begin
            regVec_318 <= _zz_regVec_0_1;
          end
          if(_zz_2[319]) begin
            regVec_319 <= _zz_regVec_0_1;
          end
          if(_zz_2[320]) begin
            regVec_320 <= _zz_regVec_0_1;
          end
          if(_zz_2[321]) begin
            regVec_321 <= _zz_regVec_0_1;
          end
          if(_zz_2[322]) begin
            regVec_322 <= _zz_regVec_0_1;
          end
          if(_zz_2[323]) begin
            regVec_323 <= _zz_regVec_0_1;
          end
          if(_zz_2[324]) begin
            regVec_324 <= _zz_regVec_0_1;
          end
          if(_zz_2[325]) begin
            regVec_325 <= _zz_regVec_0_1;
          end
          if(_zz_2[326]) begin
            regVec_326 <= _zz_regVec_0_1;
          end
          if(_zz_2[327]) begin
            regVec_327 <= _zz_regVec_0_1;
          end
          if(_zz_2[328]) begin
            regVec_328 <= _zz_regVec_0_1;
          end
          if(_zz_2[329]) begin
            regVec_329 <= _zz_regVec_0_1;
          end
          if(_zz_2[330]) begin
            regVec_330 <= _zz_regVec_0_1;
          end
          if(_zz_2[331]) begin
            regVec_331 <= _zz_regVec_0_1;
          end
          if(_zz_2[332]) begin
            regVec_332 <= _zz_regVec_0_1;
          end
          if(_zz_2[333]) begin
            regVec_333 <= _zz_regVec_0_1;
          end
          if(_zz_2[334]) begin
            regVec_334 <= _zz_regVec_0_1;
          end
          if(_zz_2[335]) begin
            regVec_335 <= _zz_regVec_0_1;
          end
          if(_zz_2[336]) begin
            regVec_336 <= _zz_regVec_0_1;
          end
          if(_zz_2[337]) begin
            regVec_337 <= _zz_regVec_0_1;
          end
          if(_zz_2[338]) begin
            regVec_338 <= _zz_regVec_0_1;
          end
          if(_zz_2[339]) begin
            regVec_339 <= _zz_regVec_0_1;
          end
          if(_zz_2[340]) begin
            regVec_340 <= _zz_regVec_0_1;
          end
          if(_zz_2[341]) begin
            regVec_341 <= _zz_regVec_0_1;
          end
          if(_zz_2[342]) begin
            regVec_342 <= _zz_regVec_0_1;
          end
          if(_zz_2[343]) begin
            regVec_343 <= _zz_regVec_0_1;
          end
          if(_zz_2[344]) begin
            regVec_344 <= _zz_regVec_0_1;
          end
          if(_zz_2[345]) begin
            regVec_345 <= _zz_regVec_0_1;
          end
          if(_zz_2[346]) begin
            regVec_346 <= _zz_regVec_0_1;
          end
          if(_zz_2[347]) begin
            regVec_347 <= _zz_regVec_0_1;
          end
          if(_zz_2[348]) begin
            regVec_348 <= _zz_regVec_0_1;
          end
          if(_zz_2[349]) begin
            regVec_349 <= _zz_regVec_0_1;
          end
          if(_zz_2[350]) begin
            regVec_350 <= _zz_regVec_0_1;
          end
          if(_zz_2[351]) begin
            regVec_351 <= _zz_regVec_0_1;
          end
          if(_zz_2[352]) begin
            regVec_352 <= _zz_regVec_0_1;
          end
          if(_zz_2[353]) begin
            regVec_353 <= _zz_regVec_0_1;
          end
          if(_zz_2[354]) begin
            regVec_354 <= _zz_regVec_0_1;
          end
          if(_zz_2[355]) begin
            regVec_355 <= _zz_regVec_0_1;
          end
          if(_zz_2[356]) begin
            regVec_356 <= _zz_regVec_0_1;
          end
          if(_zz_2[357]) begin
            regVec_357 <= _zz_regVec_0_1;
          end
          if(_zz_2[358]) begin
            regVec_358 <= _zz_regVec_0_1;
          end
          if(_zz_2[359]) begin
            regVec_359 <= _zz_regVec_0_1;
          end
          if(_zz_2[360]) begin
            regVec_360 <= _zz_regVec_0_1;
          end
          if(_zz_2[361]) begin
            regVec_361 <= _zz_regVec_0_1;
          end
          if(_zz_2[362]) begin
            regVec_362 <= _zz_regVec_0_1;
          end
          if(_zz_2[363]) begin
            regVec_363 <= _zz_regVec_0_1;
          end
          if(_zz_2[364]) begin
            regVec_364 <= _zz_regVec_0_1;
          end
          if(_zz_2[365]) begin
            regVec_365 <= _zz_regVec_0_1;
          end
          if(_zz_2[366]) begin
            regVec_366 <= _zz_regVec_0_1;
          end
          if(_zz_2[367]) begin
            regVec_367 <= _zz_regVec_0_1;
          end
          if(_zz_2[368]) begin
            regVec_368 <= _zz_regVec_0_1;
          end
          if(_zz_2[369]) begin
            regVec_369 <= _zz_regVec_0_1;
          end
          if(_zz_2[370]) begin
            regVec_370 <= _zz_regVec_0_1;
          end
          if(_zz_2[371]) begin
            regVec_371 <= _zz_regVec_0_1;
          end
          if(_zz_2[372]) begin
            regVec_372 <= _zz_regVec_0_1;
          end
          if(_zz_2[373]) begin
            regVec_373 <= _zz_regVec_0_1;
          end
          if(_zz_2[374]) begin
            regVec_374 <= _zz_regVec_0_1;
          end
          if(_zz_2[375]) begin
            regVec_375 <= _zz_regVec_0_1;
          end
          if(_zz_2[376]) begin
            regVec_376 <= _zz_regVec_0_1;
          end
          if(_zz_2[377]) begin
            regVec_377 <= _zz_regVec_0_1;
          end
          if(_zz_2[378]) begin
            regVec_378 <= _zz_regVec_0_1;
          end
          if(_zz_2[379]) begin
            regVec_379 <= _zz_regVec_0_1;
          end
          if(_zz_2[380]) begin
            regVec_380 <= _zz_regVec_0_1;
          end
          if(_zz_2[381]) begin
            regVec_381 <= _zz_regVec_0_1;
          end
          if(_zz_2[382]) begin
            regVec_382 <= _zz_regVec_0_1;
          end
          if(_zz_2[383]) begin
            regVec_383 <= _zz_regVec_0_1;
          end
          if(_zz_2[384]) begin
            regVec_384 <= _zz_regVec_0_1;
          end
          if(_zz_2[385]) begin
            regVec_385 <= _zz_regVec_0_1;
          end
          if(_zz_2[386]) begin
            regVec_386 <= _zz_regVec_0_1;
          end
          if(_zz_2[387]) begin
            regVec_387 <= _zz_regVec_0_1;
          end
          if(_zz_2[388]) begin
            regVec_388 <= _zz_regVec_0_1;
          end
          if(_zz_2[389]) begin
            regVec_389 <= _zz_regVec_0_1;
          end
          if(_zz_2[390]) begin
            regVec_390 <= _zz_regVec_0_1;
          end
          if(_zz_2[391]) begin
            regVec_391 <= _zz_regVec_0_1;
          end
          if(_zz_2[392]) begin
            regVec_392 <= _zz_regVec_0_1;
          end
          if(_zz_2[393]) begin
            regVec_393 <= _zz_regVec_0_1;
          end
          if(_zz_2[394]) begin
            regVec_394 <= _zz_regVec_0_1;
          end
          if(_zz_2[395]) begin
            regVec_395 <= _zz_regVec_0_1;
          end
          if(_zz_2[396]) begin
            regVec_396 <= _zz_regVec_0_1;
          end
          if(_zz_2[397]) begin
            regVec_397 <= _zz_regVec_0_1;
          end
          if(_zz_2[398]) begin
            regVec_398 <= _zz_regVec_0_1;
          end
          if(_zz_2[399]) begin
            regVec_399 <= _zz_regVec_0_1;
          end
          if(_zz_2[400]) begin
            regVec_400 <= _zz_regVec_0_1;
          end
          if(_zz_2[401]) begin
            regVec_401 <= _zz_regVec_0_1;
          end
          if(_zz_2[402]) begin
            regVec_402 <= _zz_regVec_0_1;
          end
          if(_zz_2[403]) begin
            regVec_403 <= _zz_regVec_0_1;
          end
          if(_zz_2[404]) begin
            regVec_404 <= _zz_regVec_0_1;
          end
          if(_zz_2[405]) begin
            regVec_405 <= _zz_regVec_0_1;
          end
          if(_zz_2[406]) begin
            regVec_406 <= _zz_regVec_0_1;
          end
          if(_zz_2[407]) begin
            regVec_407 <= _zz_regVec_0_1;
          end
          if(_zz_2[408]) begin
            regVec_408 <= _zz_regVec_0_1;
          end
          if(_zz_2[409]) begin
            regVec_409 <= _zz_regVec_0_1;
          end
          if(_zz_2[410]) begin
            regVec_410 <= _zz_regVec_0_1;
          end
          if(_zz_2[411]) begin
            regVec_411 <= _zz_regVec_0_1;
          end
          if(_zz_2[412]) begin
            regVec_412 <= _zz_regVec_0_1;
          end
          if(_zz_2[413]) begin
            regVec_413 <= _zz_regVec_0_1;
          end
          if(_zz_2[414]) begin
            regVec_414 <= _zz_regVec_0_1;
          end
          if(_zz_2[415]) begin
            regVec_415 <= _zz_regVec_0_1;
          end
          if(_zz_2[416]) begin
            regVec_416 <= _zz_regVec_0_1;
          end
          if(_zz_2[417]) begin
            regVec_417 <= _zz_regVec_0_1;
          end
          if(_zz_2[418]) begin
            regVec_418 <= _zz_regVec_0_1;
          end
          if(_zz_2[419]) begin
            regVec_419 <= _zz_regVec_0_1;
          end
          if(_zz_2[420]) begin
            regVec_420 <= _zz_regVec_0_1;
          end
          if(_zz_2[421]) begin
            regVec_421 <= _zz_regVec_0_1;
          end
          if(_zz_2[422]) begin
            regVec_422 <= _zz_regVec_0_1;
          end
          if(_zz_2[423]) begin
            regVec_423 <= _zz_regVec_0_1;
          end
          if(_zz_2[424]) begin
            regVec_424 <= _zz_regVec_0_1;
          end
          if(_zz_2[425]) begin
            regVec_425 <= _zz_regVec_0_1;
          end
          if(_zz_2[426]) begin
            regVec_426 <= _zz_regVec_0_1;
          end
          if(_zz_2[427]) begin
            regVec_427 <= _zz_regVec_0_1;
          end
          if(_zz_2[428]) begin
            regVec_428 <= _zz_regVec_0_1;
          end
          if(_zz_2[429]) begin
            regVec_429 <= _zz_regVec_0_1;
          end
          if(_zz_2[430]) begin
            regVec_430 <= _zz_regVec_0_1;
          end
          if(_zz_2[431]) begin
            regVec_431 <= _zz_regVec_0_1;
          end
          if(_zz_2[432]) begin
            regVec_432 <= _zz_regVec_0_1;
          end
          if(_zz_2[433]) begin
            regVec_433 <= _zz_regVec_0_1;
          end
          if(_zz_2[434]) begin
            regVec_434 <= _zz_regVec_0_1;
          end
          if(_zz_2[435]) begin
            regVec_435 <= _zz_regVec_0_1;
          end
          if(_zz_2[436]) begin
            regVec_436 <= _zz_regVec_0_1;
          end
          if(_zz_2[437]) begin
            regVec_437 <= _zz_regVec_0_1;
          end
          if(_zz_2[438]) begin
            regVec_438 <= _zz_regVec_0_1;
          end
          if(_zz_2[439]) begin
            regVec_439 <= _zz_regVec_0_1;
          end
          if(_zz_2[440]) begin
            regVec_440 <= _zz_regVec_0_1;
          end
          if(_zz_2[441]) begin
            regVec_441 <= _zz_regVec_0_1;
          end
          if(_zz_2[442]) begin
            regVec_442 <= _zz_regVec_0_1;
          end
          if(_zz_2[443]) begin
            regVec_443 <= _zz_regVec_0_1;
          end
          if(_zz_2[444]) begin
            regVec_444 <= _zz_regVec_0_1;
          end
          if(_zz_2[445]) begin
            regVec_445 <= _zz_regVec_0_1;
          end
          if(_zz_2[446]) begin
            regVec_446 <= _zz_regVec_0_1;
          end
          if(_zz_2[447]) begin
            regVec_447 <= _zz_regVec_0_1;
          end
          if(_zz_2[448]) begin
            regVec_448 <= _zz_regVec_0_1;
          end
          if(_zz_2[449]) begin
            regVec_449 <= _zz_regVec_0_1;
          end
          if(_zz_2[450]) begin
            regVec_450 <= _zz_regVec_0_1;
          end
          if(_zz_2[451]) begin
            regVec_451 <= _zz_regVec_0_1;
          end
          if(_zz_2[452]) begin
            regVec_452 <= _zz_regVec_0_1;
          end
          if(_zz_2[453]) begin
            regVec_453 <= _zz_regVec_0_1;
          end
          if(_zz_2[454]) begin
            regVec_454 <= _zz_regVec_0_1;
          end
          if(_zz_2[455]) begin
            regVec_455 <= _zz_regVec_0_1;
          end
          if(_zz_2[456]) begin
            regVec_456 <= _zz_regVec_0_1;
          end
          if(_zz_2[457]) begin
            regVec_457 <= _zz_regVec_0_1;
          end
          if(_zz_2[458]) begin
            regVec_458 <= _zz_regVec_0_1;
          end
          if(_zz_2[459]) begin
            regVec_459 <= _zz_regVec_0_1;
          end
          if(_zz_2[460]) begin
            regVec_460 <= _zz_regVec_0_1;
          end
          if(_zz_2[461]) begin
            regVec_461 <= _zz_regVec_0_1;
          end
          if(_zz_2[462]) begin
            regVec_462 <= _zz_regVec_0_1;
          end
          if(_zz_2[463]) begin
            regVec_463 <= _zz_regVec_0_1;
          end
          if(_zz_2[464]) begin
            regVec_464 <= _zz_regVec_0_1;
          end
          if(_zz_2[465]) begin
            regVec_465 <= _zz_regVec_0_1;
          end
          if(_zz_2[466]) begin
            regVec_466 <= _zz_regVec_0_1;
          end
          if(_zz_2[467]) begin
            regVec_467 <= _zz_regVec_0_1;
          end
          if(_zz_2[468]) begin
            regVec_468 <= _zz_regVec_0_1;
          end
          if(_zz_2[469]) begin
            regVec_469 <= _zz_regVec_0_1;
          end
          if(_zz_2[470]) begin
            regVec_470 <= _zz_regVec_0_1;
          end
          if(_zz_2[471]) begin
            regVec_471 <= _zz_regVec_0_1;
          end
          if(_zz_2[472]) begin
            regVec_472 <= _zz_regVec_0_1;
          end
          if(_zz_2[473]) begin
            regVec_473 <= _zz_regVec_0_1;
          end
          if(_zz_2[474]) begin
            regVec_474 <= _zz_regVec_0_1;
          end
          if(_zz_2[475]) begin
            regVec_475 <= _zz_regVec_0_1;
          end
          if(_zz_2[476]) begin
            regVec_476 <= _zz_regVec_0_1;
          end
          if(_zz_2[477]) begin
            regVec_477 <= _zz_regVec_0_1;
          end
          if(_zz_2[478]) begin
            regVec_478 <= _zz_regVec_0_1;
          end
          if(_zz_2[479]) begin
            regVec_479 <= _zz_regVec_0_1;
          end
          if(_zz_2[480]) begin
            regVec_480 <= _zz_regVec_0_1;
          end
          if(_zz_2[481]) begin
            regVec_481 <= _zz_regVec_0_1;
          end
          if(_zz_2[482]) begin
            regVec_482 <= _zz_regVec_0_1;
          end
          if(_zz_2[483]) begin
            regVec_483 <= _zz_regVec_0_1;
          end
          if(_zz_2[484]) begin
            regVec_484 <= _zz_regVec_0_1;
          end
          if(_zz_2[485]) begin
            regVec_485 <= _zz_regVec_0_1;
          end
          if(_zz_2[486]) begin
            regVec_486 <= _zz_regVec_0_1;
          end
          if(_zz_2[487]) begin
            regVec_487 <= _zz_regVec_0_1;
          end
          if(_zz_2[488]) begin
            regVec_488 <= _zz_regVec_0_1;
          end
          if(_zz_2[489]) begin
            regVec_489 <= _zz_regVec_0_1;
          end
          if(_zz_2[490]) begin
            regVec_490 <= _zz_regVec_0_1;
          end
          if(_zz_2[491]) begin
            regVec_491 <= _zz_regVec_0_1;
          end
          if(_zz_2[492]) begin
            regVec_492 <= _zz_regVec_0_1;
          end
          if(_zz_2[493]) begin
            regVec_493 <= _zz_regVec_0_1;
          end
          if(_zz_2[494]) begin
            regVec_494 <= _zz_regVec_0_1;
          end
          if(_zz_2[495]) begin
            regVec_495 <= _zz_regVec_0_1;
          end
          if(_zz_2[496]) begin
            regVec_496 <= _zz_regVec_0_1;
          end
          if(_zz_2[497]) begin
            regVec_497 <= _zz_regVec_0_1;
          end
          if(_zz_2[498]) begin
            regVec_498 <= _zz_regVec_0_1;
          end
          if(_zz_2[499]) begin
            regVec_499 <= _zz_regVec_0_1;
          end
          if(_zz_2[500]) begin
            regVec_500 <= _zz_regVec_0_1;
          end
          if(_zz_2[501]) begin
            regVec_501 <= _zz_regVec_0_1;
          end
          if(_zz_2[502]) begin
            regVec_502 <= _zz_regVec_0_1;
          end
          if(_zz_2[503]) begin
            regVec_503 <= _zz_regVec_0_1;
          end
          if(_zz_2[504]) begin
            regVec_504 <= _zz_regVec_0_1;
          end
          if(_zz_2[505]) begin
            regVec_505 <= _zz_regVec_0_1;
          end
          if(_zz_2[506]) begin
            regVec_506 <= _zz_regVec_0_1;
          end
          if(_zz_2[507]) begin
            regVec_507 <= _zz_regVec_0_1;
          end
          if(_zz_2[508]) begin
            regVec_508 <= _zz_regVec_0_1;
          end
          if(_zz_2[509]) begin
            regVec_509 <= _zz_regVec_0_1;
          end
          if(_zz_2[510]) begin
            regVec_510 <= _zz_regVec_0_1;
          end
          if(_zz_2[511]) begin
            regVec_511 <= _zz_regVec_0_1;
          end
          if(_zz_2[512]) begin
            regVec_512 <= _zz_regVec_0_1;
          end
          if(_zz_2[513]) begin
            regVec_513 <= _zz_regVec_0_1;
          end
          if(_zz_2[514]) begin
            regVec_514 <= _zz_regVec_0_1;
          end
          if(_zz_2[515]) begin
            regVec_515 <= _zz_regVec_0_1;
          end
          if(_zz_2[516]) begin
            regVec_516 <= _zz_regVec_0_1;
          end
          if(_zz_2[517]) begin
            regVec_517 <= _zz_regVec_0_1;
          end
          if(_zz_2[518]) begin
            regVec_518 <= _zz_regVec_0_1;
          end
          if(_zz_2[519]) begin
            regVec_519 <= _zz_regVec_0_1;
          end
          if(_zz_2[520]) begin
            regVec_520 <= _zz_regVec_0_1;
          end
          if(_zz_2[521]) begin
            regVec_521 <= _zz_regVec_0_1;
          end
          if(_zz_2[522]) begin
            regVec_522 <= _zz_regVec_0_1;
          end
          if(_zz_2[523]) begin
            regVec_523 <= _zz_regVec_0_1;
          end
          if(_zz_2[524]) begin
            regVec_524 <= _zz_regVec_0_1;
          end
          if(_zz_2[525]) begin
            regVec_525 <= _zz_regVec_0_1;
          end
          if(_zz_2[526]) begin
            regVec_526 <= _zz_regVec_0_1;
          end
          if(_zz_2[527]) begin
            regVec_527 <= _zz_regVec_0_1;
          end
          if(_zz_2[528]) begin
            regVec_528 <= _zz_regVec_0_1;
          end
          if(_zz_2[529]) begin
            regVec_529 <= _zz_regVec_0_1;
          end
          if(_zz_2[530]) begin
            regVec_530 <= _zz_regVec_0_1;
          end
          if(_zz_2[531]) begin
            regVec_531 <= _zz_regVec_0_1;
          end
          if(_zz_2[532]) begin
            regVec_532 <= _zz_regVec_0_1;
          end
          if(_zz_2[533]) begin
            regVec_533 <= _zz_regVec_0_1;
          end
          if(_zz_2[534]) begin
            regVec_534 <= _zz_regVec_0_1;
          end
          if(_zz_2[535]) begin
            regVec_535 <= _zz_regVec_0_1;
          end
          if(_zz_2[536]) begin
            regVec_536 <= _zz_regVec_0_1;
          end
          if(_zz_2[537]) begin
            regVec_537 <= _zz_regVec_0_1;
          end
          if(_zz_2[538]) begin
            regVec_538 <= _zz_regVec_0_1;
          end
          if(_zz_2[539]) begin
            regVec_539 <= _zz_regVec_0_1;
          end
          if(_zz_2[540]) begin
            regVec_540 <= _zz_regVec_0_1;
          end
          if(_zz_2[541]) begin
            regVec_541 <= _zz_regVec_0_1;
          end
          if(_zz_2[542]) begin
            regVec_542 <= _zz_regVec_0_1;
          end
          if(_zz_2[543]) begin
            regVec_543 <= _zz_regVec_0_1;
          end
          if(_zz_2[544]) begin
            regVec_544 <= _zz_regVec_0_1;
          end
          if(_zz_2[545]) begin
            regVec_545 <= _zz_regVec_0_1;
          end
          if(_zz_2[546]) begin
            regVec_546 <= _zz_regVec_0_1;
          end
          if(_zz_2[547]) begin
            regVec_547 <= _zz_regVec_0_1;
          end
          if(_zz_2[548]) begin
            regVec_548 <= _zz_regVec_0_1;
          end
          if(_zz_2[549]) begin
            regVec_549 <= _zz_regVec_0_1;
          end
          if(_zz_2[550]) begin
            regVec_550 <= _zz_regVec_0_1;
          end
          if(_zz_2[551]) begin
            regVec_551 <= _zz_regVec_0_1;
          end
          if(_zz_2[552]) begin
            regVec_552 <= _zz_regVec_0_1;
          end
          if(_zz_2[553]) begin
            regVec_553 <= _zz_regVec_0_1;
          end
          if(_zz_2[554]) begin
            regVec_554 <= _zz_regVec_0_1;
          end
          if(_zz_2[555]) begin
            regVec_555 <= _zz_regVec_0_1;
          end
          if(_zz_2[556]) begin
            regVec_556 <= _zz_regVec_0_1;
          end
          if(_zz_2[557]) begin
            regVec_557 <= _zz_regVec_0_1;
          end
          if(_zz_2[558]) begin
            regVec_558 <= _zz_regVec_0_1;
          end
          if(_zz_2[559]) begin
            regVec_559 <= _zz_regVec_0_1;
          end
          if(_zz_2[560]) begin
            regVec_560 <= _zz_regVec_0_1;
          end
          if(_zz_2[561]) begin
            regVec_561 <= _zz_regVec_0_1;
          end
          if(_zz_2[562]) begin
            regVec_562 <= _zz_regVec_0_1;
          end
          if(_zz_2[563]) begin
            regVec_563 <= _zz_regVec_0_1;
          end
          if(_zz_2[564]) begin
            regVec_564 <= _zz_regVec_0_1;
          end
          if(_zz_2[565]) begin
            regVec_565 <= _zz_regVec_0_1;
          end
          if(_zz_2[566]) begin
            regVec_566 <= _zz_regVec_0_1;
          end
          if(_zz_2[567]) begin
            regVec_567 <= _zz_regVec_0_1;
          end
          if(_zz_2[568]) begin
            regVec_568 <= _zz_regVec_0_1;
          end
          if(_zz_2[569]) begin
            regVec_569 <= _zz_regVec_0_1;
          end
          if(_zz_2[570]) begin
            regVec_570 <= _zz_regVec_0_1;
          end
          if(_zz_2[571]) begin
            regVec_571 <= _zz_regVec_0_1;
          end
          if(_zz_2[572]) begin
            regVec_572 <= _zz_regVec_0_1;
          end
          if(_zz_2[573]) begin
            regVec_573 <= _zz_regVec_0_1;
          end
          if(_zz_2[574]) begin
            regVec_574 <= _zz_regVec_0_1;
          end
          if(_zz_2[575]) begin
            regVec_575 <= _zz_regVec_0_1;
          end
          if(_zz_2[576]) begin
            regVec_576 <= _zz_regVec_0_1;
          end
          if(_zz_2[577]) begin
            regVec_577 <= _zz_regVec_0_1;
          end
          if(_zz_2[578]) begin
            regVec_578 <= _zz_regVec_0_1;
          end
          if(_zz_2[579]) begin
            regVec_579 <= _zz_regVec_0_1;
          end
          if(_zz_2[580]) begin
            regVec_580 <= _zz_regVec_0_1;
          end
          if(_zz_2[581]) begin
            regVec_581 <= _zz_regVec_0_1;
          end
          if(_zz_2[582]) begin
            regVec_582 <= _zz_regVec_0_1;
          end
          if(_zz_2[583]) begin
            regVec_583 <= _zz_regVec_0_1;
          end
          if(_zz_2[584]) begin
            regVec_584 <= _zz_regVec_0_1;
          end
          if(_zz_2[585]) begin
            regVec_585 <= _zz_regVec_0_1;
          end
          if(_zz_2[586]) begin
            regVec_586 <= _zz_regVec_0_1;
          end
          if(_zz_2[587]) begin
            regVec_587 <= _zz_regVec_0_1;
          end
          if(_zz_2[588]) begin
            regVec_588 <= _zz_regVec_0_1;
          end
          if(_zz_2[589]) begin
            regVec_589 <= _zz_regVec_0_1;
          end
          if(_zz_2[590]) begin
            regVec_590 <= _zz_regVec_0_1;
          end
          if(_zz_2[591]) begin
            regVec_591 <= _zz_regVec_0_1;
          end
          if(_zz_2[592]) begin
            regVec_592 <= _zz_regVec_0_1;
          end
          if(_zz_2[593]) begin
            regVec_593 <= _zz_regVec_0_1;
          end
          if(_zz_2[594]) begin
            regVec_594 <= _zz_regVec_0_1;
          end
          if(_zz_2[595]) begin
            regVec_595 <= _zz_regVec_0_1;
          end
          if(_zz_2[596]) begin
            regVec_596 <= _zz_regVec_0_1;
          end
          if(_zz_2[597]) begin
            regVec_597 <= _zz_regVec_0_1;
          end
          if(_zz_2[598]) begin
            regVec_598 <= _zz_regVec_0_1;
          end
          if(_zz_2[599]) begin
            regVec_599 <= _zz_regVec_0_1;
          end
          if(_zz_2[600]) begin
            regVec_600 <= _zz_regVec_0_1;
          end
          if(_zz_2[601]) begin
            regVec_601 <= _zz_regVec_0_1;
          end
          if(_zz_2[602]) begin
            regVec_602 <= _zz_regVec_0_1;
          end
          if(_zz_2[603]) begin
            regVec_603 <= _zz_regVec_0_1;
          end
          if(_zz_2[604]) begin
            regVec_604 <= _zz_regVec_0_1;
          end
          if(_zz_2[605]) begin
            regVec_605 <= _zz_regVec_0_1;
          end
          if(_zz_2[606]) begin
            regVec_606 <= _zz_regVec_0_1;
          end
          if(_zz_2[607]) begin
            regVec_607 <= _zz_regVec_0_1;
          end
          if(_zz_2[608]) begin
            regVec_608 <= _zz_regVec_0_1;
          end
          if(_zz_2[609]) begin
            regVec_609 <= _zz_regVec_0_1;
          end
          if(_zz_2[610]) begin
            regVec_610 <= _zz_regVec_0_1;
          end
          if(_zz_2[611]) begin
            regVec_611 <= _zz_regVec_0_1;
          end
          if(_zz_2[612]) begin
            regVec_612 <= _zz_regVec_0_1;
          end
          if(_zz_2[613]) begin
            regVec_613 <= _zz_regVec_0_1;
          end
          if(_zz_2[614]) begin
            regVec_614 <= _zz_regVec_0_1;
          end
          if(_zz_2[615]) begin
            regVec_615 <= _zz_regVec_0_1;
          end
          if(_zz_2[616]) begin
            regVec_616 <= _zz_regVec_0_1;
          end
          if(_zz_2[617]) begin
            regVec_617 <= _zz_regVec_0_1;
          end
          if(_zz_2[618]) begin
            regVec_618 <= _zz_regVec_0_1;
          end
          if(_zz_2[619]) begin
            regVec_619 <= _zz_regVec_0_1;
          end
          if(_zz_2[620]) begin
            regVec_620 <= _zz_regVec_0_1;
          end
          if(_zz_2[621]) begin
            regVec_621 <= _zz_regVec_0_1;
          end
          if(_zz_2[622]) begin
            regVec_622 <= _zz_regVec_0_1;
          end
          if(_zz_2[623]) begin
            regVec_623 <= _zz_regVec_0_1;
          end
          if(_zz_2[624]) begin
            regVec_624 <= _zz_regVec_0_1;
          end
          if(_zz_2[625]) begin
            regVec_625 <= _zz_regVec_0_1;
          end
          if(_zz_2[626]) begin
            regVec_626 <= _zz_regVec_0_1;
          end
          if(_zz_2[627]) begin
            regVec_627 <= _zz_regVec_0_1;
          end
          if(_zz_2[628]) begin
            regVec_628 <= _zz_regVec_0_1;
          end
          if(_zz_2[629]) begin
            regVec_629 <= _zz_regVec_0_1;
          end
          if(_zz_2[630]) begin
            regVec_630 <= _zz_regVec_0_1;
          end
          if(_zz_2[631]) begin
            regVec_631 <= _zz_regVec_0_1;
          end
          if(_zz_2[632]) begin
            regVec_632 <= _zz_regVec_0_1;
          end
          if(_zz_2[633]) begin
            regVec_633 <= _zz_regVec_0_1;
          end
          if(_zz_2[634]) begin
            regVec_634 <= _zz_regVec_0_1;
          end
          if(_zz_2[635]) begin
            regVec_635 <= _zz_regVec_0_1;
          end
          if(_zz_2[636]) begin
            regVec_636 <= _zz_regVec_0_1;
          end
          if(_zz_2[637]) begin
            regVec_637 <= _zz_regVec_0_1;
          end
          if(_zz_2[638]) begin
            regVec_638 <= _zz_regVec_0_1;
          end
          if(_zz_2[639]) begin
            regVec_639 <= _zz_regVec_0_1;
          end
          if(_zz_2[640]) begin
            regVec_640 <= _zz_regVec_0_1;
          end
          if(_zz_2[641]) begin
            regVec_641 <= _zz_regVec_0_1;
          end
          if(_zz_2[642]) begin
            regVec_642 <= _zz_regVec_0_1;
          end
          if(_zz_2[643]) begin
            regVec_643 <= _zz_regVec_0_1;
          end
          if(_zz_2[644]) begin
            regVec_644 <= _zz_regVec_0_1;
          end
          if(_zz_2[645]) begin
            regVec_645 <= _zz_regVec_0_1;
          end
          if(_zz_2[646]) begin
            regVec_646 <= _zz_regVec_0_1;
          end
          if(_zz_2[647]) begin
            regVec_647 <= _zz_regVec_0_1;
          end
          if(_zz_2[648]) begin
            regVec_648 <= _zz_regVec_0_1;
          end
          if(_zz_2[649]) begin
            regVec_649 <= _zz_regVec_0_1;
          end
          if(_zz_2[650]) begin
            regVec_650 <= _zz_regVec_0_1;
          end
          if(_zz_2[651]) begin
            regVec_651 <= _zz_regVec_0_1;
          end
          if(_zz_2[652]) begin
            regVec_652 <= _zz_regVec_0_1;
          end
          if(_zz_2[653]) begin
            regVec_653 <= _zz_regVec_0_1;
          end
          if(_zz_2[654]) begin
            regVec_654 <= _zz_regVec_0_1;
          end
          if(_zz_2[655]) begin
            regVec_655 <= _zz_regVec_0_1;
          end
          if(_zz_2[656]) begin
            regVec_656 <= _zz_regVec_0_1;
          end
          if(_zz_2[657]) begin
            regVec_657 <= _zz_regVec_0_1;
          end
          if(_zz_2[658]) begin
            regVec_658 <= _zz_regVec_0_1;
          end
          if(_zz_2[659]) begin
            regVec_659 <= _zz_regVec_0_1;
          end
          if(_zz_2[660]) begin
            regVec_660 <= _zz_regVec_0_1;
          end
          if(_zz_2[661]) begin
            regVec_661 <= _zz_regVec_0_1;
          end
          if(_zz_2[662]) begin
            regVec_662 <= _zz_regVec_0_1;
          end
          if(_zz_2[663]) begin
            regVec_663 <= _zz_regVec_0_1;
          end
          if(_zz_2[664]) begin
            regVec_664 <= _zz_regVec_0_1;
          end
          if(_zz_2[665]) begin
            regVec_665 <= _zz_regVec_0_1;
          end
          if(_zz_2[666]) begin
            regVec_666 <= _zz_regVec_0_1;
          end
          if(_zz_2[667]) begin
            regVec_667 <= _zz_regVec_0_1;
          end
          if(_zz_2[668]) begin
            regVec_668 <= _zz_regVec_0_1;
          end
          if(_zz_2[669]) begin
            regVec_669 <= _zz_regVec_0_1;
          end
          if(_zz_2[670]) begin
            regVec_670 <= _zz_regVec_0_1;
          end
          if(_zz_2[671]) begin
            regVec_671 <= _zz_regVec_0_1;
          end
          if(_zz_2[672]) begin
            regVec_672 <= _zz_regVec_0_1;
          end
          if(_zz_2[673]) begin
            regVec_673 <= _zz_regVec_0_1;
          end
          if(_zz_2[674]) begin
            regVec_674 <= _zz_regVec_0_1;
          end
          if(_zz_2[675]) begin
            regVec_675 <= _zz_regVec_0_1;
          end
          if(_zz_2[676]) begin
            regVec_676 <= _zz_regVec_0_1;
          end
          if(_zz_2[677]) begin
            regVec_677 <= _zz_regVec_0_1;
          end
          if(_zz_2[678]) begin
            regVec_678 <= _zz_regVec_0_1;
          end
          if(_zz_2[679]) begin
            regVec_679 <= _zz_regVec_0_1;
          end
          if(_zz_2[680]) begin
            regVec_680 <= _zz_regVec_0_1;
          end
          if(_zz_2[681]) begin
            regVec_681 <= _zz_regVec_0_1;
          end
          if(_zz_2[682]) begin
            regVec_682 <= _zz_regVec_0_1;
          end
          if(_zz_2[683]) begin
            regVec_683 <= _zz_regVec_0_1;
          end
          if(_zz_2[684]) begin
            regVec_684 <= _zz_regVec_0_1;
          end
          if(_zz_2[685]) begin
            regVec_685 <= _zz_regVec_0_1;
          end
          if(_zz_2[686]) begin
            regVec_686 <= _zz_regVec_0_1;
          end
          if(_zz_2[687]) begin
            regVec_687 <= _zz_regVec_0_1;
          end
          if(_zz_2[688]) begin
            regVec_688 <= _zz_regVec_0_1;
          end
          if(_zz_2[689]) begin
            regVec_689 <= _zz_regVec_0_1;
          end
          if(_zz_2[690]) begin
            regVec_690 <= _zz_regVec_0_1;
          end
          if(_zz_2[691]) begin
            regVec_691 <= _zz_regVec_0_1;
          end
          if(_zz_2[692]) begin
            regVec_692 <= _zz_regVec_0_1;
          end
          if(_zz_2[693]) begin
            regVec_693 <= _zz_regVec_0_1;
          end
          if(_zz_2[694]) begin
            regVec_694 <= _zz_regVec_0_1;
          end
          if(_zz_2[695]) begin
            regVec_695 <= _zz_regVec_0_1;
          end
          if(_zz_2[696]) begin
            regVec_696 <= _zz_regVec_0_1;
          end
          if(_zz_2[697]) begin
            regVec_697 <= _zz_regVec_0_1;
          end
          if(_zz_2[698]) begin
            regVec_698 <= _zz_regVec_0_1;
          end
          if(_zz_2[699]) begin
            regVec_699 <= _zz_regVec_0_1;
          end
          if(_zz_2[700]) begin
            regVec_700 <= _zz_regVec_0_1;
          end
          if(_zz_2[701]) begin
            regVec_701 <= _zz_regVec_0_1;
          end
          if(_zz_2[702]) begin
            regVec_702 <= _zz_regVec_0_1;
          end
          if(_zz_2[703]) begin
            regVec_703 <= _zz_regVec_0_1;
          end
          if(_zz_2[704]) begin
            regVec_704 <= _zz_regVec_0_1;
          end
          if(_zz_2[705]) begin
            regVec_705 <= _zz_regVec_0_1;
          end
          if(_zz_2[706]) begin
            regVec_706 <= _zz_regVec_0_1;
          end
          if(_zz_2[707]) begin
            regVec_707 <= _zz_regVec_0_1;
          end
          if(_zz_2[708]) begin
            regVec_708 <= _zz_regVec_0_1;
          end
          if(_zz_2[709]) begin
            regVec_709 <= _zz_regVec_0_1;
          end
          if(_zz_2[710]) begin
            regVec_710 <= _zz_regVec_0_1;
          end
          if(_zz_2[711]) begin
            regVec_711 <= _zz_regVec_0_1;
          end
          if(_zz_2[712]) begin
            regVec_712 <= _zz_regVec_0_1;
          end
          if(_zz_2[713]) begin
            regVec_713 <= _zz_regVec_0_1;
          end
          if(_zz_2[714]) begin
            regVec_714 <= _zz_regVec_0_1;
          end
          if(_zz_2[715]) begin
            regVec_715 <= _zz_regVec_0_1;
          end
          if(_zz_2[716]) begin
            regVec_716 <= _zz_regVec_0_1;
          end
          if(_zz_2[717]) begin
            regVec_717 <= _zz_regVec_0_1;
          end
          if(_zz_2[718]) begin
            regVec_718 <= _zz_regVec_0_1;
          end
          if(_zz_2[719]) begin
            regVec_719 <= _zz_regVec_0_1;
          end
          if(_zz_2[720]) begin
            regVec_720 <= _zz_regVec_0_1;
          end
          if(_zz_2[721]) begin
            regVec_721 <= _zz_regVec_0_1;
          end
          if(_zz_2[722]) begin
            regVec_722 <= _zz_regVec_0_1;
          end
          if(_zz_2[723]) begin
            regVec_723 <= _zz_regVec_0_1;
          end
          if(_zz_2[724]) begin
            regVec_724 <= _zz_regVec_0_1;
          end
          if(_zz_2[725]) begin
            regVec_725 <= _zz_regVec_0_1;
          end
          if(_zz_2[726]) begin
            regVec_726 <= _zz_regVec_0_1;
          end
          if(_zz_2[727]) begin
            regVec_727 <= _zz_regVec_0_1;
          end
          if(_zz_2[728]) begin
            regVec_728 <= _zz_regVec_0_1;
          end
          if(_zz_2[729]) begin
            regVec_729 <= _zz_regVec_0_1;
          end
          if(_zz_2[730]) begin
            regVec_730 <= _zz_regVec_0_1;
          end
          if(_zz_2[731]) begin
            regVec_731 <= _zz_regVec_0_1;
          end
          if(_zz_2[732]) begin
            regVec_732 <= _zz_regVec_0_1;
          end
          if(_zz_2[733]) begin
            regVec_733 <= _zz_regVec_0_1;
          end
          if(_zz_2[734]) begin
            regVec_734 <= _zz_regVec_0_1;
          end
          if(_zz_2[735]) begin
            regVec_735 <= _zz_regVec_0_1;
          end
          if(_zz_2[736]) begin
            regVec_736 <= _zz_regVec_0_1;
          end
          if(_zz_2[737]) begin
            regVec_737 <= _zz_regVec_0_1;
          end
          if(_zz_2[738]) begin
            regVec_738 <= _zz_regVec_0_1;
          end
          if(_zz_2[739]) begin
            regVec_739 <= _zz_regVec_0_1;
          end
          if(_zz_2[740]) begin
            regVec_740 <= _zz_regVec_0_1;
          end
          if(_zz_2[741]) begin
            regVec_741 <= _zz_regVec_0_1;
          end
          if(_zz_2[742]) begin
            regVec_742 <= _zz_regVec_0_1;
          end
          if(_zz_2[743]) begin
            regVec_743 <= _zz_regVec_0_1;
          end
          if(_zz_2[744]) begin
            regVec_744 <= _zz_regVec_0_1;
          end
          if(_zz_2[745]) begin
            regVec_745 <= _zz_regVec_0_1;
          end
          if(_zz_2[746]) begin
            regVec_746 <= _zz_regVec_0_1;
          end
          if(_zz_2[747]) begin
            regVec_747 <= _zz_regVec_0_1;
          end
          if(_zz_2[748]) begin
            regVec_748 <= _zz_regVec_0_1;
          end
          if(_zz_2[749]) begin
            regVec_749 <= _zz_regVec_0_1;
          end
          if(_zz_2[750]) begin
            regVec_750 <= _zz_regVec_0_1;
          end
          if(_zz_2[751]) begin
            regVec_751 <= _zz_regVec_0_1;
          end
          if(_zz_2[752]) begin
            regVec_752 <= _zz_regVec_0_1;
          end
          if(_zz_2[753]) begin
            regVec_753 <= _zz_regVec_0_1;
          end
          if(_zz_2[754]) begin
            regVec_754 <= _zz_regVec_0_1;
          end
          if(_zz_2[755]) begin
            regVec_755 <= _zz_regVec_0_1;
          end
          if(_zz_2[756]) begin
            regVec_756 <= _zz_regVec_0_1;
          end
          if(_zz_2[757]) begin
            regVec_757 <= _zz_regVec_0_1;
          end
          if(_zz_2[758]) begin
            regVec_758 <= _zz_regVec_0_1;
          end
          if(_zz_2[759]) begin
            regVec_759 <= _zz_regVec_0_1;
          end
          if(_zz_2[760]) begin
            regVec_760 <= _zz_regVec_0_1;
          end
          if(_zz_2[761]) begin
            regVec_761 <= _zz_regVec_0_1;
          end
          if(_zz_2[762]) begin
            regVec_762 <= _zz_regVec_0_1;
          end
          if(_zz_2[763]) begin
            regVec_763 <= _zz_regVec_0_1;
          end
          if(_zz_2[764]) begin
            regVec_764 <= _zz_regVec_0_1;
          end
          if(_zz_2[765]) begin
            regVec_765 <= _zz_regVec_0_1;
          end
          if(_zz_2[766]) begin
            regVec_766 <= _zz_regVec_0_1;
          end
          if(_zz_2[767]) begin
            regVec_767 <= _zz_regVec_0_1;
          end
          if(_zz_2[768]) begin
            regVec_768 <= _zz_regVec_0_1;
          end
          if(_zz_2[769]) begin
            regVec_769 <= _zz_regVec_0_1;
          end
          if(_zz_2[770]) begin
            regVec_770 <= _zz_regVec_0_1;
          end
          if(_zz_2[771]) begin
            regVec_771 <= _zz_regVec_0_1;
          end
          if(_zz_2[772]) begin
            regVec_772 <= _zz_regVec_0_1;
          end
          if(_zz_2[773]) begin
            regVec_773 <= _zz_regVec_0_1;
          end
          if(_zz_2[774]) begin
            regVec_774 <= _zz_regVec_0_1;
          end
          if(_zz_2[775]) begin
            regVec_775 <= _zz_regVec_0_1;
          end
          if(_zz_2[776]) begin
            regVec_776 <= _zz_regVec_0_1;
          end
          if(_zz_2[777]) begin
            regVec_777 <= _zz_regVec_0_1;
          end
          if(_zz_2[778]) begin
            regVec_778 <= _zz_regVec_0_1;
          end
          if(_zz_2[779]) begin
            regVec_779 <= _zz_regVec_0_1;
          end
          if(_zz_2[780]) begin
            regVec_780 <= _zz_regVec_0_1;
          end
          if(_zz_2[781]) begin
            regVec_781 <= _zz_regVec_0_1;
          end
          if(_zz_2[782]) begin
            regVec_782 <= _zz_regVec_0_1;
          end
          if(_zz_2[783]) begin
            regVec_783 <= _zz_regVec_0_1;
          end
          if(_zz_2[784]) begin
            regVec_784 <= _zz_regVec_0_1;
          end
          if(_zz_2[785]) begin
            regVec_785 <= _zz_regVec_0_1;
          end
          if(_zz_2[786]) begin
            regVec_786 <= _zz_regVec_0_1;
          end
          if(_zz_2[787]) begin
            regVec_787 <= _zz_regVec_0_1;
          end
          if(_zz_2[788]) begin
            regVec_788 <= _zz_regVec_0_1;
          end
          if(_zz_2[789]) begin
            regVec_789 <= _zz_regVec_0_1;
          end
          if(_zz_2[790]) begin
            regVec_790 <= _zz_regVec_0_1;
          end
          if(_zz_2[791]) begin
            regVec_791 <= _zz_regVec_0_1;
          end
          if(_zz_2[792]) begin
            regVec_792 <= _zz_regVec_0_1;
          end
          if(_zz_2[793]) begin
            regVec_793 <= _zz_regVec_0_1;
          end
          if(_zz_2[794]) begin
            regVec_794 <= _zz_regVec_0_1;
          end
          if(_zz_2[795]) begin
            regVec_795 <= _zz_regVec_0_1;
          end
          if(_zz_2[796]) begin
            regVec_796 <= _zz_regVec_0_1;
          end
          if(_zz_2[797]) begin
            regVec_797 <= _zz_regVec_0_1;
          end
          if(_zz_2[798]) begin
            regVec_798 <= _zz_regVec_0_1;
          end
          if(_zz_2[799]) begin
            regVec_799 <= _zz_regVec_0_1;
          end
          if(_zz_2[800]) begin
            regVec_800 <= _zz_regVec_0_1;
          end
          if(_zz_2[801]) begin
            regVec_801 <= _zz_regVec_0_1;
          end
          if(_zz_2[802]) begin
            regVec_802 <= _zz_regVec_0_1;
          end
          if(_zz_2[803]) begin
            regVec_803 <= _zz_regVec_0_1;
          end
          if(_zz_2[804]) begin
            regVec_804 <= _zz_regVec_0_1;
          end
          if(_zz_2[805]) begin
            regVec_805 <= _zz_regVec_0_1;
          end
          if(_zz_2[806]) begin
            regVec_806 <= _zz_regVec_0_1;
          end
          if(_zz_2[807]) begin
            regVec_807 <= _zz_regVec_0_1;
          end
          if(_zz_2[808]) begin
            regVec_808 <= _zz_regVec_0_1;
          end
          if(_zz_2[809]) begin
            regVec_809 <= _zz_regVec_0_1;
          end
          if(_zz_2[810]) begin
            regVec_810 <= _zz_regVec_0_1;
          end
          if(_zz_2[811]) begin
            regVec_811 <= _zz_regVec_0_1;
          end
          if(_zz_2[812]) begin
            regVec_812 <= _zz_regVec_0_1;
          end
          if(_zz_2[813]) begin
            regVec_813 <= _zz_regVec_0_1;
          end
          if(_zz_2[814]) begin
            regVec_814 <= _zz_regVec_0_1;
          end
          if(_zz_2[815]) begin
            regVec_815 <= _zz_regVec_0_1;
          end
          if(_zz_2[816]) begin
            regVec_816 <= _zz_regVec_0_1;
          end
          if(_zz_2[817]) begin
            regVec_817 <= _zz_regVec_0_1;
          end
          if(_zz_2[818]) begin
            regVec_818 <= _zz_regVec_0_1;
          end
          if(_zz_2[819]) begin
            regVec_819 <= _zz_regVec_0_1;
          end
          if(_zz_2[820]) begin
            regVec_820 <= _zz_regVec_0_1;
          end
          if(_zz_2[821]) begin
            regVec_821 <= _zz_regVec_0_1;
          end
          if(_zz_2[822]) begin
            regVec_822 <= _zz_regVec_0_1;
          end
          if(_zz_2[823]) begin
            regVec_823 <= _zz_regVec_0_1;
          end
          if(_zz_2[824]) begin
            regVec_824 <= _zz_regVec_0_1;
          end
          if(_zz_2[825]) begin
            regVec_825 <= _zz_regVec_0_1;
          end
          if(_zz_2[826]) begin
            regVec_826 <= _zz_regVec_0_1;
          end
          if(_zz_2[827]) begin
            regVec_827 <= _zz_regVec_0_1;
          end
          if(_zz_2[828]) begin
            regVec_828 <= _zz_regVec_0_1;
          end
          if(_zz_2[829]) begin
            regVec_829 <= _zz_regVec_0_1;
          end
          if(_zz_2[830]) begin
            regVec_830 <= _zz_regVec_0_1;
          end
          if(_zz_2[831]) begin
            regVec_831 <= _zz_regVec_0_1;
          end
          if(_zz_2[832]) begin
            regVec_832 <= _zz_regVec_0_1;
          end
          if(_zz_2[833]) begin
            regVec_833 <= _zz_regVec_0_1;
          end
          if(_zz_2[834]) begin
            regVec_834 <= _zz_regVec_0_1;
          end
          if(_zz_2[835]) begin
            regVec_835 <= _zz_regVec_0_1;
          end
          if(_zz_2[836]) begin
            regVec_836 <= _zz_regVec_0_1;
          end
          if(_zz_2[837]) begin
            regVec_837 <= _zz_regVec_0_1;
          end
          if(_zz_2[838]) begin
            regVec_838 <= _zz_regVec_0_1;
          end
          if(_zz_2[839]) begin
            regVec_839 <= _zz_regVec_0_1;
          end
          if(_zz_2[840]) begin
            regVec_840 <= _zz_regVec_0_1;
          end
          if(_zz_2[841]) begin
            regVec_841 <= _zz_regVec_0_1;
          end
          if(_zz_2[842]) begin
            regVec_842 <= _zz_regVec_0_1;
          end
          if(_zz_2[843]) begin
            regVec_843 <= _zz_regVec_0_1;
          end
          if(_zz_2[844]) begin
            regVec_844 <= _zz_regVec_0_1;
          end
          if(_zz_2[845]) begin
            regVec_845 <= _zz_regVec_0_1;
          end
          if(_zz_2[846]) begin
            regVec_846 <= _zz_regVec_0_1;
          end
          if(_zz_2[847]) begin
            regVec_847 <= _zz_regVec_0_1;
          end
          if(_zz_2[848]) begin
            regVec_848 <= _zz_regVec_0_1;
          end
          if(_zz_2[849]) begin
            regVec_849 <= _zz_regVec_0_1;
          end
          if(_zz_2[850]) begin
            regVec_850 <= _zz_regVec_0_1;
          end
          if(_zz_2[851]) begin
            regVec_851 <= _zz_regVec_0_1;
          end
          if(_zz_2[852]) begin
            regVec_852 <= _zz_regVec_0_1;
          end
          if(_zz_2[853]) begin
            regVec_853 <= _zz_regVec_0_1;
          end
          if(_zz_2[854]) begin
            regVec_854 <= _zz_regVec_0_1;
          end
          if(_zz_2[855]) begin
            regVec_855 <= _zz_regVec_0_1;
          end
          if(_zz_2[856]) begin
            regVec_856 <= _zz_regVec_0_1;
          end
          if(_zz_2[857]) begin
            regVec_857 <= _zz_regVec_0_1;
          end
          if(_zz_2[858]) begin
            regVec_858 <= _zz_regVec_0_1;
          end
          if(_zz_2[859]) begin
            regVec_859 <= _zz_regVec_0_1;
          end
          if(_zz_2[860]) begin
            regVec_860 <= _zz_regVec_0_1;
          end
          if(_zz_2[861]) begin
            regVec_861 <= _zz_regVec_0_1;
          end
          if(_zz_2[862]) begin
            regVec_862 <= _zz_regVec_0_1;
          end
          if(_zz_2[863]) begin
            regVec_863 <= _zz_regVec_0_1;
          end
          if(_zz_2[864]) begin
            regVec_864 <= _zz_regVec_0_1;
          end
          if(_zz_2[865]) begin
            regVec_865 <= _zz_regVec_0_1;
          end
          if(_zz_2[866]) begin
            regVec_866 <= _zz_regVec_0_1;
          end
          if(_zz_2[867]) begin
            regVec_867 <= _zz_regVec_0_1;
          end
          if(_zz_2[868]) begin
            regVec_868 <= _zz_regVec_0_1;
          end
          if(_zz_2[869]) begin
            regVec_869 <= _zz_regVec_0_1;
          end
          if(_zz_2[870]) begin
            regVec_870 <= _zz_regVec_0_1;
          end
          if(_zz_2[871]) begin
            regVec_871 <= _zz_regVec_0_1;
          end
          if(_zz_2[872]) begin
            regVec_872 <= _zz_regVec_0_1;
          end
          if(_zz_2[873]) begin
            regVec_873 <= _zz_regVec_0_1;
          end
          if(_zz_2[874]) begin
            regVec_874 <= _zz_regVec_0_1;
          end
          if(_zz_2[875]) begin
            regVec_875 <= _zz_regVec_0_1;
          end
          if(_zz_2[876]) begin
            regVec_876 <= _zz_regVec_0_1;
          end
          if(_zz_2[877]) begin
            regVec_877 <= _zz_regVec_0_1;
          end
          if(_zz_2[878]) begin
            regVec_878 <= _zz_regVec_0_1;
          end
          if(_zz_2[879]) begin
            regVec_879 <= _zz_regVec_0_1;
          end
          if(_zz_2[880]) begin
            regVec_880 <= _zz_regVec_0_1;
          end
          if(_zz_2[881]) begin
            regVec_881 <= _zz_regVec_0_1;
          end
          if(_zz_2[882]) begin
            regVec_882 <= _zz_regVec_0_1;
          end
          if(_zz_2[883]) begin
            regVec_883 <= _zz_regVec_0_1;
          end
          if(_zz_2[884]) begin
            regVec_884 <= _zz_regVec_0_1;
          end
          if(_zz_2[885]) begin
            regVec_885 <= _zz_regVec_0_1;
          end
          if(_zz_2[886]) begin
            regVec_886 <= _zz_regVec_0_1;
          end
          if(_zz_2[887]) begin
            regVec_887 <= _zz_regVec_0_1;
          end
          if(_zz_2[888]) begin
            regVec_888 <= _zz_regVec_0_1;
          end
          if(_zz_2[889]) begin
            regVec_889 <= _zz_regVec_0_1;
          end
          if(_zz_2[890]) begin
            regVec_890 <= _zz_regVec_0_1;
          end
          if(_zz_2[891]) begin
            regVec_891 <= _zz_regVec_0_1;
          end
          if(_zz_2[892]) begin
            regVec_892 <= _zz_regVec_0_1;
          end
          if(_zz_2[893]) begin
            regVec_893 <= _zz_regVec_0_1;
          end
          if(_zz_2[894]) begin
            regVec_894 <= _zz_regVec_0_1;
          end
          if(_zz_2[895]) begin
            regVec_895 <= _zz_regVec_0_1;
          end
          if(_zz_2[896]) begin
            regVec_896 <= _zz_regVec_0_1;
          end
          if(_zz_2[897]) begin
            regVec_897 <= _zz_regVec_0_1;
          end
          if(_zz_2[898]) begin
            regVec_898 <= _zz_regVec_0_1;
          end
          if(_zz_2[899]) begin
            regVec_899 <= _zz_regVec_0_1;
          end
          if(_zz_2[900]) begin
            regVec_900 <= _zz_regVec_0_1;
          end
          if(_zz_2[901]) begin
            regVec_901 <= _zz_regVec_0_1;
          end
          if(_zz_2[902]) begin
            regVec_902 <= _zz_regVec_0_1;
          end
          if(_zz_2[903]) begin
            regVec_903 <= _zz_regVec_0_1;
          end
          if(_zz_2[904]) begin
            regVec_904 <= _zz_regVec_0_1;
          end
          if(_zz_2[905]) begin
            regVec_905 <= _zz_regVec_0_1;
          end
          if(_zz_2[906]) begin
            regVec_906 <= _zz_regVec_0_1;
          end
          if(_zz_2[907]) begin
            regVec_907 <= _zz_regVec_0_1;
          end
          if(_zz_2[908]) begin
            regVec_908 <= _zz_regVec_0_1;
          end
          if(_zz_2[909]) begin
            regVec_909 <= _zz_regVec_0_1;
          end
          if(_zz_2[910]) begin
            regVec_910 <= _zz_regVec_0_1;
          end
          if(_zz_2[911]) begin
            regVec_911 <= _zz_regVec_0_1;
          end
          if(_zz_2[912]) begin
            regVec_912 <= _zz_regVec_0_1;
          end
          if(_zz_2[913]) begin
            regVec_913 <= _zz_regVec_0_1;
          end
          if(_zz_2[914]) begin
            regVec_914 <= _zz_regVec_0_1;
          end
          if(_zz_2[915]) begin
            regVec_915 <= _zz_regVec_0_1;
          end
          if(_zz_2[916]) begin
            regVec_916 <= _zz_regVec_0_1;
          end
          if(_zz_2[917]) begin
            regVec_917 <= _zz_regVec_0_1;
          end
          if(_zz_2[918]) begin
            regVec_918 <= _zz_regVec_0_1;
          end
          if(_zz_2[919]) begin
            regVec_919 <= _zz_regVec_0_1;
          end
          if(_zz_2[920]) begin
            regVec_920 <= _zz_regVec_0_1;
          end
          if(_zz_2[921]) begin
            regVec_921 <= _zz_regVec_0_1;
          end
          if(_zz_2[922]) begin
            regVec_922 <= _zz_regVec_0_1;
          end
          if(_zz_2[923]) begin
            regVec_923 <= _zz_regVec_0_1;
          end
          if(_zz_2[924]) begin
            regVec_924 <= _zz_regVec_0_1;
          end
          if(_zz_2[925]) begin
            regVec_925 <= _zz_regVec_0_1;
          end
          if(_zz_2[926]) begin
            regVec_926 <= _zz_regVec_0_1;
          end
          if(_zz_2[927]) begin
            regVec_927 <= _zz_regVec_0_1;
          end
          if(_zz_2[928]) begin
            regVec_928 <= _zz_regVec_0_1;
          end
          if(_zz_2[929]) begin
            regVec_929 <= _zz_regVec_0_1;
          end
          if(_zz_2[930]) begin
            regVec_930 <= _zz_regVec_0_1;
          end
          if(_zz_2[931]) begin
            regVec_931 <= _zz_regVec_0_1;
          end
          if(_zz_2[932]) begin
            regVec_932 <= _zz_regVec_0_1;
          end
          if(_zz_2[933]) begin
            regVec_933 <= _zz_regVec_0_1;
          end
          if(_zz_2[934]) begin
            regVec_934 <= _zz_regVec_0_1;
          end
          if(_zz_2[935]) begin
            regVec_935 <= _zz_regVec_0_1;
          end
          if(_zz_2[936]) begin
            regVec_936 <= _zz_regVec_0_1;
          end
          if(_zz_2[937]) begin
            regVec_937 <= _zz_regVec_0_1;
          end
          if(_zz_2[938]) begin
            regVec_938 <= _zz_regVec_0_1;
          end
          if(_zz_2[939]) begin
            regVec_939 <= _zz_regVec_0_1;
          end
          if(_zz_2[940]) begin
            regVec_940 <= _zz_regVec_0_1;
          end
          if(_zz_2[941]) begin
            regVec_941 <= _zz_regVec_0_1;
          end
          if(_zz_2[942]) begin
            regVec_942 <= _zz_regVec_0_1;
          end
          if(_zz_2[943]) begin
            regVec_943 <= _zz_regVec_0_1;
          end
          if(_zz_2[944]) begin
            regVec_944 <= _zz_regVec_0_1;
          end
          if(_zz_2[945]) begin
            regVec_945 <= _zz_regVec_0_1;
          end
          if(_zz_2[946]) begin
            regVec_946 <= _zz_regVec_0_1;
          end
          if(_zz_2[947]) begin
            regVec_947 <= _zz_regVec_0_1;
          end
          if(_zz_2[948]) begin
            regVec_948 <= _zz_regVec_0_1;
          end
          if(_zz_2[949]) begin
            regVec_949 <= _zz_regVec_0_1;
          end
          if(_zz_2[950]) begin
            regVec_950 <= _zz_regVec_0_1;
          end
          if(_zz_2[951]) begin
            regVec_951 <= _zz_regVec_0_1;
          end
          if(_zz_2[952]) begin
            regVec_952 <= _zz_regVec_0_1;
          end
          if(_zz_2[953]) begin
            regVec_953 <= _zz_regVec_0_1;
          end
          if(_zz_2[954]) begin
            regVec_954 <= _zz_regVec_0_1;
          end
          if(_zz_2[955]) begin
            regVec_955 <= _zz_regVec_0_1;
          end
          if(_zz_2[956]) begin
            regVec_956 <= _zz_regVec_0_1;
          end
          if(_zz_2[957]) begin
            regVec_957 <= _zz_regVec_0_1;
          end
          if(_zz_2[958]) begin
            regVec_958 <= _zz_regVec_0_1;
          end
          if(_zz_2[959]) begin
            regVec_959 <= _zz_regVec_0_1;
          end
          if(_zz_2[960]) begin
            regVec_960 <= _zz_regVec_0_1;
          end
          if(_zz_2[961]) begin
            regVec_961 <= _zz_regVec_0_1;
          end
          if(_zz_2[962]) begin
            regVec_962 <= _zz_regVec_0_1;
          end
          if(_zz_2[963]) begin
            regVec_963 <= _zz_regVec_0_1;
          end
          if(_zz_2[964]) begin
            regVec_964 <= _zz_regVec_0_1;
          end
          if(_zz_2[965]) begin
            regVec_965 <= _zz_regVec_0_1;
          end
          if(_zz_2[966]) begin
            regVec_966 <= _zz_regVec_0_1;
          end
          if(_zz_2[967]) begin
            regVec_967 <= _zz_regVec_0_1;
          end
          if(_zz_2[968]) begin
            regVec_968 <= _zz_regVec_0_1;
          end
          if(_zz_2[969]) begin
            regVec_969 <= _zz_regVec_0_1;
          end
          if(_zz_2[970]) begin
            regVec_970 <= _zz_regVec_0_1;
          end
          if(_zz_2[971]) begin
            regVec_971 <= _zz_regVec_0_1;
          end
          if(_zz_2[972]) begin
            regVec_972 <= _zz_regVec_0_1;
          end
          if(_zz_2[973]) begin
            regVec_973 <= _zz_regVec_0_1;
          end
          if(_zz_2[974]) begin
            regVec_974 <= _zz_regVec_0_1;
          end
          if(_zz_2[975]) begin
            regVec_975 <= _zz_regVec_0_1;
          end
          if(_zz_2[976]) begin
            regVec_976 <= _zz_regVec_0_1;
          end
          if(_zz_2[977]) begin
            regVec_977 <= _zz_regVec_0_1;
          end
          if(_zz_2[978]) begin
            regVec_978 <= _zz_regVec_0_1;
          end
          if(_zz_2[979]) begin
            regVec_979 <= _zz_regVec_0_1;
          end
          if(_zz_2[980]) begin
            regVec_980 <= _zz_regVec_0_1;
          end
          if(_zz_2[981]) begin
            regVec_981 <= _zz_regVec_0_1;
          end
          if(_zz_2[982]) begin
            regVec_982 <= _zz_regVec_0_1;
          end
          if(_zz_2[983]) begin
            regVec_983 <= _zz_regVec_0_1;
          end
          if(_zz_2[984]) begin
            regVec_984 <= _zz_regVec_0_1;
          end
          if(_zz_2[985]) begin
            regVec_985 <= _zz_regVec_0_1;
          end
          if(_zz_2[986]) begin
            regVec_986 <= _zz_regVec_0_1;
          end
          if(_zz_2[987]) begin
            regVec_987 <= _zz_regVec_0_1;
          end
          if(_zz_2[988]) begin
            regVec_988 <= _zz_regVec_0_1;
          end
          if(_zz_2[989]) begin
            regVec_989 <= _zz_regVec_0_1;
          end
          if(_zz_2[990]) begin
            regVec_990 <= _zz_regVec_0_1;
          end
          if(_zz_2[991]) begin
            regVec_991 <= _zz_regVec_0_1;
          end
          if(_zz_2[992]) begin
            regVec_992 <= _zz_regVec_0_1;
          end
          if(_zz_2[993]) begin
            regVec_993 <= _zz_regVec_0_1;
          end
          if(_zz_2[994]) begin
            regVec_994 <= _zz_regVec_0_1;
          end
          if(_zz_2[995]) begin
            regVec_995 <= _zz_regVec_0_1;
          end
          if(_zz_2[996]) begin
            regVec_996 <= _zz_regVec_0_1;
          end
          if(_zz_2[997]) begin
            regVec_997 <= _zz_regVec_0_1;
          end
          if(_zz_2[998]) begin
            regVec_998 <= _zz_regVec_0_1;
          end
          if(_zz_2[999]) begin
            regVec_999 <= _zz_regVec_0_1;
          end
          if(_zz_2[1000]) begin
            regVec_1000 <= _zz_regVec_0_1;
          end
          if(_zz_2[1001]) begin
            regVec_1001 <= _zz_regVec_0_1;
          end
          if(_zz_2[1002]) begin
            regVec_1002 <= _zz_regVec_0_1;
          end
          if(_zz_2[1003]) begin
            regVec_1003 <= _zz_regVec_0_1;
          end
          if(_zz_2[1004]) begin
            regVec_1004 <= _zz_regVec_0_1;
          end
          if(_zz_2[1005]) begin
            regVec_1005 <= _zz_regVec_0_1;
          end
          if(_zz_2[1006]) begin
            regVec_1006 <= _zz_regVec_0_1;
          end
          if(_zz_2[1007]) begin
            regVec_1007 <= _zz_regVec_0_1;
          end
          if(_zz_2[1008]) begin
            regVec_1008 <= _zz_regVec_0_1;
          end
          if(_zz_2[1009]) begin
            regVec_1009 <= _zz_regVec_0_1;
          end
          if(_zz_2[1010]) begin
            regVec_1010 <= _zz_regVec_0_1;
          end
          if(_zz_2[1011]) begin
            regVec_1011 <= _zz_regVec_0_1;
          end
          if(_zz_2[1012]) begin
            regVec_1012 <= _zz_regVec_0_1;
          end
          if(_zz_2[1013]) begin
            regVec_1013 <= _zz_regVec_0_1;
          end
          if(_zz_2[1014]) begin
            regVec_1014 <= _zz_regVec_0_1;
          end
          if(_zz_2[1015]) begin
            regVec_1015 <= _zz_regVec_0_1;
          end
          if(_zz_2[1016]) begin
            regVec_1016 <= _zz_regVec_0_1;
          end
          if(_zz_2[1017]) begin
            regVec_1017 <= _zz_regVec_0_1;
          end
          if(_zz_2[1018]) begin
            regVec_1018 <= _zz_regVec_0_1;
          end
          if(_zz_2[1019]) begin
            regVec_1019 <= _zz_regVec_0_1;
          end
          if(_zz_2[1020]) begin
            regVec_1020 <= _zz_regVec_0_1;
          end
          if(_zz_2[1021]) begin
            regVec_1021 <= _zz_regVec_0_1;
          end
          if(_zz_2[1022]) begin
            regVec_1022 <= _zz_regVec_0_1;
          end
          if(_zz_2[1023]) begin
            regVec_1023 <= _zz_regVec_0_1;
          end
          if(_zz_2[1024]) begin
            regVec_1024 <= _zz_regVec_0_1;
          end
          if(_zz_2[1025]) begin
            regVec_1025 <= _zz_regVec_0_1;
          end
          if(_zz_2[1026]) begin
            regVec_1026 <= _zz_regVec_0_1;
          end
          if(_zz_2[1027]) begin
            regVec_1027 <= _zz_regVec_0_1;
          end
          if(_zz_2[1028]) begin
            regVec_1028 <= _zz_regVec_0_1;
          end
          if(_zz_2[1029]) begin
            regVec_1029 <= _zz_regVec_0_1;
          end
          if(_zz_2[1030]) begin
            regVec_1030 <= _zz_regVec_0_1;
          end
          if(_zz_2[1031]) begin
            regVec_1031 <= _zz_regVec_0_1;
          end
          if(_zz_2[1032]) begin
            regVec_1032 <= _zz_regVec_0_1;
          end
          if(_zz_2[1033]) begin
            regVec_1033 <= _zz_regVec_0_1;
          end
          if(_zz_2[1034]) begin
            regVec_1034 <= _zz_regVec_0_1;
          end
          if(_zz_2[1035]) begin
            regVec_1035 <= _zz_regVec_0_1;
          end
          if(_zz_2[1036]) begin
            regVec_1036 <= _zz_regVec_0_1;
          end
          if(_zz_2[1037]) begin
            regVec_1037 <= _zz_regVec_0_1;
          end
          if(_zz_2[1038]) begin
            regVec_1038 <= _zz_regVec_0_1;
          end
          if(_zz_2[1039]) begin
            regVec_1039 <= _zz_regVec_0_1;
          end
          if(_zz_2[1040]) begin
            regVec_1040 <= _zz_regVec_0_1;
          end
          if(_zz_2[1041]) begin
            regVec_1041 <= _zz_regVec_0_1;
          end
          if(_zz_2[1042]) begin
            regVec_1042 <= _zz_regVec_0_1;
          end
          if(_zz_2[1043]) begin
            regVec_1043 <= _zz_regVec_0_1;
          end
          if(_zz_2[1044]) begin
            regVec_1044 <= _zz_regVec_0_1;
          end
          if(_zz_2[1045]) begin
            regVec_1045 <= _zz_regVec_0_1;
          end
          if(_zz_2[1046]) begin
            regVec_1046 <= _zz_regVec_0_1;
          end
          if(_zz_2[1047]) begin
            regVec_1047 <= _zz_regVec_0_1;
          end
          if(_zz_2[1048]) begin
            regVec_1048 <= _zz_regVec_0_1;
          end
          if(_zz_2[1049]) begin
            regVec_1049 <= _zz_regVec_0_1;
          end
          if(_zz_2[1050]) begin
            regVec_1050 <= _zz_regVec_0_1;
          end
          if(_zz_2[1051]) begin
            regVec_1051 <= _zz_regVec_0_1;
          end
          if(_zz_2[1052]) begin
            regVec_1052 <= _zz_regVec_0_1;
          end
          if(_zz_2[1053]) begin
            regVec_1053 <= _zz_regVec_0_1;
          end
          if(_zz_2[1054]) begin
            regVec_1054 <= _zz_regVec_0_1;
          end
          if(_zz_2[1055]) begin
            regVec_1055 <= _zz_regVec_0_1;
          end
          if(_zz_2[1056]) begin
            regVec_1056 <= _zz_regVec_0_1;
          end
          if(_zz_2[1057]) begin
            regVec_1057 <= _zz_regVec_0_1;
          end
          if(_zz_2[1058]) begin
            regVec_1058 <= _zz_regVec_0_1;
          end
          if(_zz_2[1059]) begin
            regVec_1059 <= _zz_regVec_0_1;
          end
          if(_zz_2[1060]) begin
            regVec_1060 <= _zz_regVec_0_1;
          end
          if(_zz_2[1061]) begin
            regVec_1061 <= _zz_regVec_0_1;
          end
          if(_zz_2[1062]) begin
            regVec_1062 <= _zz_regVec_0_1;
          end
          if(_zz_2[1063]) begin
            regVec_1063 <= _zz_regVec_0_1;
          end
          if(_zz_2[1064]) begin
            regVec_1064 <= _zz_regVec_0_1;
          end
          if(_zz_2[1065]) begin
            regVec_1065 <= _zz_regVec_0_1;
          end
          if(_zz_2[1066]) begin
            regVec_1066 <= _zz_regVec_0_1;
          end
          if(_zz_2[1067]) begin
            regVec_1067 <= _zz_regVec_0_1;
          end
          if(_zz_2[1068]) begin
            regVec_1068 <= _zz_regVec_0_1;
          end
          if(_zz_2[1069]) begin
            regVec_1069 <= _zz_regVec_0_1;
          end
          if(_zz_2[1070]) begin
            regVec_1070 <= _zz_regVec_0_1;
          end
          if(_zz_2[1071]) begin
            regVec_1071 <= _zz_regVec_0_1;
          end
          if(_zz_2[1072]) begin
            regVec_1072 <= _zz_regVec_0_1;
          end
          if(_zz_2[1073]) begin
            regVec_1073 <= _zz_regVec_0_1;
          end
          if(_zz_2[1074]) begin
            regVec_1074 <= _zz_regVec_0_1;
          end
          if(_zz_2[1075]) begin
            regVec_1075 <= _zz_regVec_0_1;
          end
          if(_zz_2[1076]) begin
            regVec_1076 <= _zz_regVec_0_1;
          end
          if(_zz_2[1077]) begin
            regVec_1077 <= _zz_regVec_0_1;
          end
          if(_zz_2[1078]) begin
            regVec_1078 <= _zz_regVec_0_1;
          end
          if(_zz_2[1079]) begin
            regVec_1079 <= _zz_regVec_0_1;
          end
          if(_zz_2[1080]) begin
            regVec_1080 <= _zz_regVec_0_1;
          end
          if(_zz_2[1081]) begin
            regVec_1081 <= _zz_regVec_0_1;
          end
          if(_zz_2[1082]) begin
            regVec_1082 <= _zz_regVec_0_1;
          end
          if(_zz_2[1083]) begin
            regVec_1083 <= _zz_regVec_0_1;
          end
          if(_zz_2[1084]) begin
            regVec_1084 <= _zz_regVec_0_1;
          end
          if(_zz_2[1085]) begin
            regVec_1085 <= _zz_regVec_0_1;
          end
          if(_zz_2[1086]) begin
            regVec_1086 <= _zz_regVec_0_1;
          end
          if(_zz_2[1087]) begin
            regVec_1087 <= _zz_regVec_0_1;
          end
          if(_zz_2[1088]) begin
            regVec_1088 <= _zz_regVec_0_1;
          end
          if(_zz_2[1089]) begin
            regVec_1089 <= _zz_regVec_0_1;
          end
          if(_zz_2[1090]) begin
            regVec_1090 <= _zz_regVec_0_1;
          end
          if(_zz_2[1091]) begin
            regVec_1091 <= _zz_regVec_0_1;
          end
          if(_zz_2[1092]) begin
            regVec_1092 <= _zz_regVec_0_1;
          end
          if(_zz_2[1093]) begin
            regVec_1093 <= _zz_regVec_0_1;
          end
          if(_zz_2[1094]) begin
            regVec_1094 <= _zz_regVec_0_1;
          end
          if(_zz_2[1095]) begin
            regVec_1095 <= _zz_regVec_0_1;
          end
          if(_zz_2[1096]) begin
            regVec_1096 <= _zz_regVec_0_1;
          end
          if(_zz_2[1097]) begin
            regVec_1097 <= _zz_regVec_0_1;
          end
          if(_zz_2[1098]) begin
            regVec_1098 <= _zz_regVec_0_1;
          end
          if(_zz_2[1099]) begin
            regVec_1099 <= _zz_regVec_0_1;
          end
          if(_zz_2[1100]) begin
            regVec_1100 <= _zz_regVec_0_1;
          end
          if(_zz_2[1101]) begin
            regVec_1101 <= _zz_regVec_0_1;
          end
          if(_zz_2[1102]) begin
            regVec_1102 <= _zz_regVec_0_1;
          end
          if(_zz_2[1103]) begin
            regVec_1103 <= _zz_regVec_0_1;
          end
          if(_zz_2[1104]) begin
            regVec_1104 <= _zz_regVec_0_1;
          end
          if(_zz_2[1105]) begin
            regVec_1105 <= _zz_regVec_0_1;
          end
          if(_zz_2[1106]) begin
            regVec_1106 <= _zz_regVec_0_1;
          end
          if(_zz_2[1107]) begin
            regVec_1107 <= _zz_regVec_0_1;
          end
          if(_zz_2[1108]) begin
            regVec_1108 <= _zz_regVec_0_1;
          end
          if(_zz_2[1109]) begin
            regVec_1109 <= _zz_regVec_0_1;
          end
          if(_zz_2[1110]) begin
            regVec_1110 <= _zz_regVec_0_1;
          end
          if(_zz_2[1111]) begin
            regVec_1111 <= _zz_regVec_0_1;
          end
          if(_zz_2[1112]) begin
            regVec_1112 <= _zz_regVec_0_1;
          end
          if(_zz_2[1113]) begin
            regVec_1113 <= _zz_regVec_0_1;
          end
          if(_zz_2[1114]) begin
            regVec_1114 <= _zz_regVec_0_1;
          end
          if(_zz_2[1115]) begin
            regVec_1115 <= _zz_regVec_0_1;
          end
          if(_zz_2[1116]) begin
            regVec_1116 <= _zz_regVec_0_1;
          end
          if(_zz_2[1117]) begin
            regVec_1117 <= _zz_regVec_0_1;
          end
          if(_zz_2[1118]) begin
            regVec_1118 <= _zz_regVec_0_1;
          end
          if(_zz_2[1119]) begin
            regVec_1119 <= _zz_regVec_0_1;
          end
          if(_zz_2[1120]) begin
            regVec_1120 <= _zz_regVec_0_1;
          end
          if(_zz_2[1121]) begin
            regVec_1121 <= _zz_regVec_0_1;
          end
          if(_zz_2[1122]) begin
            regVec_1122 <= _zz_regVec_0_1;
          end
          if(_zz_2[1123]) begin
            regVec_1123 <= _zz_regVec_0_1;
          end
          if(_zz_2[1124]) begin
            regVec_1124 <= _zz_regVec_0_1;
          end
          if(_zz_2[1125]) begin
            regVec_1125 <= _zz_regVec_0_1;
          end
          if(_zz_2[1126]) begin
            regVec_1126 <= _zz_regVec_0_1;
          end
          if(_zz_2[1127]) begin
            regVec_1127 <= _zz_regVec_0_1;
          end
          if(_zz_2[1128]) begin
            regVec_1128 <= _zz_regVec_0_1;
          end
          if(_zz_2[1129]) begin
            regVec_1129 <= _zz_regVec_0_1;
          end
          if(_zz_2[1130]) begin
            regVec_1130 <= _zz_regVec_0_1;
          end
          if(_zz_2[1131]) begin
            regVec_1131 <= _zz_regVec_0_1;
          end
          if(_zz_2[1132]) begin
            regVec_1132 <= _zz_regVec_0_1;
          end
          if(_zz_2[1133]) begin
            regVec_1133 <= _zz_regVec_0_1;
          end
          if(_zz_2[1134]) begin
            regVec_1134 <= _zz_regVec_0_1;
          end
          if(_zz_2[1135]) begin
            regVec_1135 <= _zz_regVec_0_1;
          end
          if(_zz_2[1136]) begin
            regVec_1136 <= _zz_regVec_0_1;
          end
          if(_zz_2[1137]) begin
            regVec_1137 <= _zz_regVec_0_1;
          end
          if(_zz_2[1138]) begin
            regVec_1138 <= _zz_regVec_0_1;
          end
          if(_zz_2[1139]) begin
            regVec_1139 <= _zz_regVec_0_1;
          end
          if(_zz_2[1140]) begin
            regVec_1140 <= _zz_regVec_0_1;
          end
          if(_zz_2[1141]) begin
            regVec_1141 <= _zz_regVec_0_1;
          end
          if(_zz_2[1142]) begin
            regVec_1142 <= _zz_regVec_0_1;
          end
          if(_zz_2[1143]) begin
            regVec_1143 <= _zz_regVec_0_1;
          end
          if(_zz_2[1144]) begin
            regVec_1144 <= _zz_regVec_0_1;
          end
          if(_zz_2[1145]) begin
            regVec_1145 <= _zz_regVec_0_1;
          end
          if(_zz_2[1146]) begin
            regVec_1146 <= _zz_regVec_0_1;
          end
          if(_zz_2[1147]) begin
            regVec_1147 <= _zz_regVec_0_1;
          end
          if(_zz_2[1148]) begin
            regVec_1148 <= _zz_regVec_0_1;
          end
          if(_zz_2[1149]) begin
            regVec_1149 <= _zz_regVec_0_1;
          end
          if(_zz_2[1150]) begin
            regVec_1150 <= _zz_regVec_0_1;
          end
          if(_zz_2[1151]) begin
            regVec_1151 <= _zz_regVec_0_1;
          end
          if(_zz_2[1152]) begin
            regVec_1152 <= _zz_regVec_0_1;
          end
          if(_zz_2[1153]) begin
            regVec_1153 <= _zz_regVec_0_1;
          end
          if(_zz_2[1154]) begin
            regVec_1154 <= _zz_regVec_0_1;
          end
          if(_zz_2[1155]) begin
            regVec_1155 <= _zz_regVec_0_1;
          end
          if(_zz_2[1156]) begin
            regVec_1156 <= _zz_regVec_0_1;
          end
          if(_zz_2[1157]) begin
            regVec_1157 <= _zz_regVec_0_1;
          end
          if(_zz_2[1158]) begin
            regVec_1158 <= _zz_regVec_0_1;
          end
          if(_zz_2[1159]) begin
            regVec_1159 <= _zz_regVec_0_1;
          end
          if(_zz_2[1160]) begin
            regVec_1160 <= _zz_regVec_0_1;
          end
          if(_zz_2[1161]) begin
            regVec_1161 <= _zz_regVec_0_1;
          end
          if(_zz_2[1162]) begin
            regVec_1162 <= _zz_regVec_0_1;
          end
          if(_zz_2[1163]) begin
            regVec_1163 <= _zz_regVec_0_1;
          end
          if(_zz_2[1164]) begin
            regVec_1164 <= _zz_regVec_0_1;
          end
          if(_zz_2[1165]) begin
            regVec_1165 <= _zz_regVec_0_1;
          end
          if(_zz_2[1166]) begin
            regVec_1166 <= _zz_regVec_0_1;
          end
          if(_zz_2[1167]) begin
            regVec_1167 <= _zz_regVec_0_1;
          end
          if(_zz_2[1168]) begin
            regVec_1168 <= _zz_regVec_0_1;
          end
          if(_zz_2[1169]) begin
            regVec_1169 <= _zz_regVec_0_1;
          end
          if(_zz_2[1170]) begin
            regVec_1170 <= _zz_regVec_0_1;
          end
          if(_zz_2[1171]) begin
            regVec_1171 <= _zz_regVec_0_1;
          end
          if(_zz_2[1172]) begin
            regVec_1172 <= _zz_regVec_0_1;
          end
          if(_zz_2[1173]) begin
            regVec_1173 <= _zz_regVec_0_1;
          end
          if(_zz_2[1174]) begin
            regVec_1174 <= _zz_regVec_0_1;
          end
          if(_zz_2[1175]) begin
            regVec_1175 <= _zz_regVec_0_1;
          end
          if(_zz_2[1176]) begin
            regVec_1176 <= _zz_regVec_0_1;
          end
          if(_zz_2[1177]) begin
            regVec_1177 <= _zz_regVec_0_1;
          end
          if(_zz_2[1178]) begin
            regVec_1178 <= _zz_regVec_0_1;
          end
          if(_zz_2[1179]) begin
            regVec_1179 <= _zz_regVec_0_1;
          end
          if(_zz_2[1180]) begin
            regVec_1180 <= _zz_regVec_0_1;
          end
          if(_zz_2[1181]) begin
            regVec_1181 <= _zz_regVec_0_1;
          end
          if(_zz_2[1182]) begin
            regVec_1182 <= _zz_regVec_0_1;
          end
          if(_zz_2[1183]) begin
            regVec_1183 <= _zz_regVec_0_1;
          end
          if(_zz_2[1184]) begin
            regVec_1184 <= _zz_regVec_0_1;
          end
          if(_zz_2[1185]) begin
            regVec_1185 <= _zz_regVec_0_1;
          end
          if(_zz_2[1186]) begin
            regVec_1186 <= _zz_regVec_0_1;
          end
          if(_zz_2[1187]) begin
            regVec_1187 <= _zz_regVec_0_1;
          end
          if(_zz_2[1188]) begin
            regVec_1188 <= _zz_regVec_0_1;
          end
          if(_zz_2[1189]) begin
            regVec_1189 <= _zz_regVec_0_1;
          end
          if(_zz_2[1190]) begin
            regVec_1190 <= _zz_regVec_0_1;
          end
          if(_zz_2[1191]) begin
            regVec_1191 <= _zz_regVec_0_1;
          end
          if(_zz_2[1192]) begin
            regVec_1192 <= _zz_regVec_0_1;
          end
          if(_zz_2[1193]) begin
            regVec_1193 <= _zz_regVec_0_1;
          end
          if(_zz_2[1194]) begin
            regVec_1194 <= _zz_regVec_0_1;
          end
          if(_zz_2[1195]) begin
            regVec_1195 <= _zz_regVec_0_1;
          end
          if(_zz_2[1196]) begin
            regVec_1196 <= _zz_regVec_0_1;
          end
          if(_zz_2[1197]) begin
            regVec_1197 <= _zz_regVec_0_1;
          end
          if(_zz_2[1198]) begin
            regVec_1198 <= _zz_regVec_0_1;
          end
          if(_zz_2[1199]) begin
            regVec_1199 <= _zz_regVec_0_1;
          end
          if(_zz_2[1200]) begin
            regVec_1200 <= _zz_regVec_0_1;
          end
          if(_zz_2[1201]) begin
            regVec_1201 <= _zz_regVec_0_1;
          end
          if(_zz_2[1202]) begin
            regVec_1202 <= _zz_regVec_0_1;
          end
          if(_zz_2[1203]) begin
            regVec_1203 <= _zz_regVec_0_1;
          end
          if(_zz_2[1204]) begin
            regVec_1204 <= _zz_regVec_0_1;
          end
          if(_zz_2[1205]) begin
            regVec_1205 <= _zz_regVec_0_1;
          end
          if(_zz_2[1206]) begin
            regVec_1206 <= _zz_regVec_0_1;
          end
          if(_zz_2[1207]) begin
            regVec_1207 <= _zz_regVec_0_1;
          end
          if(_zz_2[1208]) begin
            regVec_1208 <= _zz_regVec_0_1;
          end
          if(_zz_2[1209]) begin
            regVec_1209 <= _zz_regVec_0_1;
          end
          if(_zz_2[1210]) begin
            regVec_1210 <= _zz_regVec_0_1;
          end
          if(_zz_2[1211]) begin
            regVec_1211 <= _zz_regVec_0_1;
          end
          if(_zz_2[1212]) begin
            regVec_1212 <= _zz_regVec_0_1;
          end
          if(_zz_2[1213]) begin
            regVec_1213 <= _zz_regVec_0_1;
          end
          if(_zz_2[1214]) begin
            regVec_1214 <= _zz_regVec_0_1;
          end
          if(_zz_2[1215]) begin
            regVec_1215 <= _zz_regVec_0_1;
          end
          if(_zz_2[1216]) begin
            regVec_1216 <= _zz_regVec_0_1;
          end
          if(_zz_2[1217]) begin
            regVec_1217 <= _zz_regVec_0_1;
          end
          if(_zz_2[1218]) begin
            regVec_1218 <= _zz_regVec_0_1;
          end
          if(_zz_2[1219]) begin
            regVec_1219 <= _zz_regVec_0_1;
          end
          if(_zz_2[1220]) begin
            regVec_1220 <= _zz_regVec_0_1;
          end
          if(_zz_2[1221]) begin
            regVec_1221 <= _zz_regVec_0_1;
          end
          if(_zz_2[1222]) begin
            regVec_1222 <= _zz_regVec_0_1;
          end
          if(_zz_2[1223]) begin
            regVec_1223 <= _zz_regVec_0_1;
          end
          if(_zz_2[1224]) begin
            regVec_1224 <= _zz_regVec_0_1;
          end
          if(_zz_2[1225]) begin
            regVec_1225 <= _zz_regVec_0_1;
          end
          if(_zz_2[1226]) begin
            regVec_1226 <= _zz_regVec_0_1;
          end
          if(_zz_2[1227]) begin
            regVec_1227 <= _zz_regVec_0_1;
          end
          if(_zz_2[1228]) begin
            regVec_1228 <= _zz_regVec_0_1;
          end
          if(_zz_2[1229]) begin
            regVec_1229 <= _zz_regVec_0_1;
          end
          if(_zz_2[1230]) begin
            regVec_1230 <= _zz_regVec_0_1;
          end
          if(_zz_2[1231]) begin
            regVec_1231 <= _zz_regVec_0_1;
          end
          if(_zz_2[1232]) begin
            regVec_1232 <= _zz_regVec_0_1;
          end
          if(_zz_2[1233]) begin
            regVec_1233 <= _zz_regVec_0_1;
          end
          if(_zz_2[1234]) begin
            regVec_1234 <= _zz_regVec_0_1;
          end
          if(_zz_2[1235]) begin
            regVec_1235 <= _zz_regVec_0_1;
          end
          if(_zz_2[1236]) begin
            regVec_1236 <= _zz_regVec_0_1;
          end
          if(_zz_2[1237]) begin
            regVec_1237 <= _zz_regVec_0_1;
          end
          if(_zz_2[1238]) begin
            regVec_1238 <= _zz_regVec_0_1;
          end
          if(_zz_2[1239]) begin
            regVec_1239 <= _zz_regVec_0_1;
          end
          if(_zz_2[1240]) begin
            regVec_1240 <= _zz_regVec_0_1;
          end
          if(_zz_2[1241]) begin
            regVec_1241 <= _zz_regVec_0_1;
          end
          if(_zz_2[1242]) begin
            regVec_1242 <= _zz_regVec_0_1;
          end
          if(_zz_2[1243]) begin
            regVec_1243 <= _zz_regVec_0_1;
          end
          if(_zz_2[1244]) begin
            regVec_1244 <= _zz_regVec_0_1;
          end
          if(_zz_2[1245]) begin
            regVec_1245 <= _zz_regVec_0_1;
          end
          if(_zz_2[1246]) begin
            regVec_1246 <= _zz_regVec_0_1;
          end
          if(_zz_2[1247]) begin
            regVec_1247 <= _zz_regVec_0_1;
          end
          if(_zz_2[1248]) begin
            regVec_1248 <= _zz_regVec_0_1;
          end
          if(_zz_2[1249]) begin
            regVec_1249 <= _zz_regVec_0_1;
          end
          if(_zz_2[1250]) begin
            regVec_1250 <= _zz_regVec_0_1;
          end
          if(_zz_2[1251]) begin
            regVec_1251 <= _zz_regVec_0_1;
          end
          if(_zz_2[1252]) begin
            regVec_1252 <= _zz_regVec_0_1;
          end
          if(_zz_2[1253]) begin
            regVec_1253 <= _zz_regVec_0_1;
          end
          if(_zz_2[1254]) begin
            regVec_1254 <= _zz_regVec_0_1;
          end
          if(_zz_2[1255]) begin
            regVec_1255 <= _zz_regVec_0_1;
          end
          if(_zz_2[1256]) begin
            regVec_1256 <= _zz_regVec_0_1;
          end
          if(_zz_2[1257]) begin
            regVec_1257 <= _zz_regVec_0_1;
          end
          if(_zz_2[1258]) begin
            regVec_1258 <= _zz_regVec_0_1;
          end
          if(_zz_2[1259]) begin
            regVec_1259 <= _zz_regVec_0_1;
          end
          if(_zz_2[1260]) begin
            regVec_1260 <= _zz_regVec_0_1;
          end
          if(_zz_2[1261]) begin
            regVec_1261 <= _zz_regVec_0_1;
          end
          if(_zz_2[1262]) begin
            regVec_1262 <= _zz_regVec_0_1;
          end
          if(_zz_2[1263]) begin
            regVec_1263 <= _zz_regVec_0_1;
          end
          if(_zz_2[1264]) begin
            regVec_1264 <= _zz_regVec_0_1;
          end
          if(_zz_2[1265]) begin
            regVec_1265 <= _zz_regVec_0_1;
          end
          if(_zz_2[1266]) begin
            regVec_1266 <= _zz_regVec_0_1;
          end
          if(_zz_2[1267]) begin
            regVec_1267 <= _zz_regVec_0_1;
          end
          if(_zz_2[1268]) begin
            regVec_1268 <= _zz_regVec_0_1;
          end
          if(_zz_2[1269]) begin
            regVec_1269 <= _zz_regVec_0_1;
          end
          if(_zz_2[1270]) begin
            regVec_1270 <= _zz_regVec_0_1;
          end
          if(_zz_2[1271]) begin
            regVec_1271 <= _zz_regVec_0_1;
          end
          if(_zz_2[1272]) begin
            regVec_1272 <= _zz_regVec_0_1;
          end
          if(_zz_2[1273]) begin
            regVec_1273 <= _zz_regVec_0_1;
          end
          if(_zz_2[1274]) begin
            regVec_1274 <= _zz_regVec_0_1;
          end
          if(_zz_2[1275]) begin
            regVec_1275 <= _zz_regVec_0_1;
          end
          if(_zz_2[1276]) begin
            regVec_1276 <= _zz_regVec_0_1;
          end
          if(_zz_2[1277]) begin
            regVec_1277 <= _zz_regVec_0_1;
          end
          if(_zz_2[1278]) begin
            regVec_1278 <= _zz_regVec_0_1;
          end
          if(_zz_2[1279]) begin
            regVec_1279 <= _zz_regVec_0_1;
          end
          if(_zz_2[1280]) begin
            regVec_1280 <= _zz_regVec_0_1;
          end
          if(_zz_2[1281]) begin
            regVec_1281 <= _zz_regVec_0_1;
          end
          if(_zz_2[1282]) begin
            regVec_1282 <= _zz_regVec_0_1;
          end
          if(_zz_2[1283]) begin
            regVec_1283 <= _zz_regVec_0_1;
          end
          if(_zz_2[1284]) begin
            regVec_1284 <= _zz_regVec_0_1;
          end
          if(_zz_2[1285]) begin
            regVec_1285 <= _zz_regVec_0_1;
          end
          if(_zz_2[1286]) begin
            regVec_1286 <= _zz_regVec_0_1;
          end
          if(_zz_2[1287]) begin
            regVec_1287 <= _zz_regVec_0_1;
          end
          if(_zz_2[1288]) begin
            regVec_1288 <= _zz_regVec_0_1;
          end
          if(_zz_2[1289]) begin
            regVec_1289 <= _zz_regVec_0_1;
          end
          if(_zz_2[1290]) begin
            regVec_1290 <= _zz_regVec_0_1;
          end
          if(_zz_2[1291]) begin
            regVec_1291 <= _zz_regVec_0_1;
          end
          if(_zz_2[1292]) begin
            regVec_1292 <= _zz_regVec_0_1;
          end
          if(_zz_2[1293]) begin
            regVec_1293 <= _zz_regVec_0_1;
          end
          if(_zz_2[1294]) begin
            regVec_1294 <= _zz_regVec_0_1;
          end
          if(_zz_2[1295]) begin
            regVec_1295 <= _zz_regVec_0_1;
          end
          if(_zz_2[1296]) begin
            regVec_1296 <= _zz_regVec_0_1;
          end
          if(_zz_2[1297]) begin
            regVec_1297 <= _zz_regVec_0_1;
          end
          if(_zz_2[1298]) begin
            regVec_1298 <= _zz_regVec_0_1;
          end
          if(_zz_2[1299]) begin
            regVec_1299 <= _zz_regVec_0_1;
          end
          if(_zz_2[1300]) begin
            regVec_1300 <= _zz_regVec_0_1;
          end
          if(_zz_2[1301]) begin
            regVec_1301 <= _zz_regVec_0_1;
          end
          if(_zz_2[1302]) begin
            regVec_1302 <= _zz_regVec_0_1;
          end
          if(_zz_2[1303]) begin
            regVec_1303 <= _zz_regVec_0_1;
          end
          if(_zz_2[1304]) begin
            regVec_1304 <= _zz_regVec_0_1;
          end
          if(_zz_2[1305]) begin
            regVec_1305 <= _zz_regVec_0_1;
          end
          if(_zz_2[1306]) begin
            regVec_1306 <= _zz_regVec_0_1;
          end
          if(_zz_2[1307]) begin
            regVec_1307 <= _zz_regVec_0_1;
          end
          if(_zz_2[1308]) begin
            regVec_1308 <= _zz_regVec_0_1;
          end
          if(_zz_2[1309]) begin
            regVec_1309 <= _zz_regVec_0_1;
          end
          if(_zz_2[1310]) begin
            regVec_1310 <= _zz_regVec_0_1;
          end
          if(_zz_2[1311]) begin
            regVec_1311 <= _zz_regVec_0_1;
          end
          if(_zz_2[1312]) begin
            regVec_1312 <= _zz_regVec_0_1;
          end
          if(_zz_2[1313]) begin
            regVec_1313 <= _zz_regVec_0_1;
          end
          if(_zz_2[1314]) begin
            regVec_1314 <= _zz_regVec_0_1;
          end
          if(_zz_2[1315]) begin
            regVec_1315 <= _zz_regVec_0_1;
          end
          if(_zz_2[1316]) begin
            regVec_1316 <= _zz_regVec_0_1;
          end
          if(_zz_2[1317]) begin
            regVec_1317 <= _zz_regVec_0_1;
          end
          if(_zz_2[1318]) begin
            regVec_1318 <= _zz_regVec_0_1;
          end
          if(_zz_2[1319]) begin
            regVec_1319 <= _zz_regVec_0_1;
          end
          if(_zz_2[1320]) begin
            regVec_1320 <= _zz_regVec_0_1;
          end
          if(_zz_2[1321]) begin
            regVec_1321 <= _zz_regVec_0_1;
          end
          if(_zz_2[1322]) begin
            regVec_1322 <= _zz_regVec_0_1;
          end
          if(_zz_2[1323]) begin
            regVec_1323 <= _zz_regVec_0_1;
          end
          if(_zz_2[1324]) begin
            regVec_1324 <= _zz_regVec_0_1;
          end
          if(_zz_2[1325]) begin
            regVec_1325 <= _zz_regVec_0_1;
          end
          if(_zz_2[1326]) begin
            regVec_1326 <= _zz_regVec_0_1;
          end
          if(_zz_2[1327]) begin
            regVec_1327 <= _zz_regVec_0_1;
          end
          if(_zz_2[1328]) begin
            regVec_1328 <= _zz_regVec_0_1;
          end
          if(_zz_2[1329]) begin
            regVec_1329 <= _zz_regVec_0_1;
          end
          if(_zz_2[1330]) begin
            regVec_1330 <= _zz_regVec_0_1;
          end
          if(_zz_2[1331]) begin
            regVec_1331 <= _zz_regVec_0_1;
          end
          if(_zz_2[1332]) begin
            regVec_1332 <= _zz_regVec_0_1;
          end
          if(_zz_2[1333]) begin
            regVec_1333 <= _zz_regVec_0_1;
          end
          if(_zz_2[1334]) begin
            regVec_1334 <= _zz_regVec_0_1;
          end
          if(_zz_2[1335]) begin
            regVec_1335 <= _zz_regVec_0_1;
          end
          if(_zz_2[1336]) begin
            regVec_1336 <= _zz_regVec_0_1;
          end
          if(_zz_2[1337]) begin
            regVec_1337 <= _zz_regVec_0_1;
          end
          if(_zz_2[1338]) begin
            regVec_1338 <= _zz_regVec_0_1;
          end
          if(_zz_2[1339]) begin
            regVec_1339 <= _zz_regVec_0_1;
          end
          if(_zz_2[1340]) begin
            regVec_1340 <= _zz_regVec_0_1;
          end
          if(_zz_2[1341]) begin
            regVec_1341 <= _zz_regVec_0_1;
          end
          if(_zz_2[1342]) begin
            regVec_1342 <= _zz_regVec_0_1;
          end
          if(_zz_2[1343]) begin
            regVec_1343 <= _zz_regVec_0_1;
          end
          if(_zz_2[1344]) begin
            regVec_1344 <= _zz_regVec_0_1;
          end
          if(_zz_2[1345]) begin
            regVec_1345 <= _zz_regVec_0_1;
          end
          if(_zz_2[1346]) begin
            regVec_1346 <= _zz_regVec_0_1;
          end
          if(_zz_2[1347]) begin
            regVec_1347 <= _zz_regVec_0_1;
          end
          if(_zz_2[1348]) begin
            regVec_1348 <= _zz_regVec_0_1;
          end
          if(_zz_2[1349]) begin
            regVec_1349 <= _zz_regVec_0_1;
          end
          if(_zz_2[1350]) begin
            regVec_1350 <= _zz_regVec_0_1;
          end
          if(_zz_2[1351]) begin
            regVec_1351 <= _zz_regVec_0_1;
          end
          if(_zz_2[1352]) begin
            regVec_1352 <= _zz_regVec_0_1;
          end
          if(_zz_2[1353]) begin
            regVec_1353 <= _zz_regVec_0_1;
          end
          if(_zz_2[1354]) begin
            regVec_1354 <= _zz_regVec_0_1;
          end
          if(_zz_2[1355]) begin
            regVec_1355 <= _zz_regVec_0_1;
          end
          if(_zz_2[1356]) begin
            regVec_1356 <= _zz_regVec_0_1;
          end
          if(_zz_2[1357]) begin
            regVec_1357 <= _zz_regVec_0_1;
          end
          if(_zz_2[1358]) begin
            regVec_1358 <= _zz_regVec_0_1;
          end
          if(_zz_2[1359]) begin
            regVec_1359 <= _zz_regVec_0_1;
          end
          if(_zz_2[1360]) begin
            regVec_1360 <= _zz_regVec_0_1;
          end
          if(_zz_2[1361]) begin
            regVec_1361 <= _zz_regVec_0_1;
          end
          if(_zz_2[1362]) begin
            regVec_1362 <= _zz_regVec_0_1;
          end
          if(_zz_2[1363]) begin
            regVec_1363 <= _zz_regVec_0_1;
          end
          if(_zz_2[1364]) begin
            regVec_1364 <= _zz_regVec_0_1;
          end
          if(_zz_2[1365]) begin
            regVec_1365 <= _zz_regVec_0_1;
          end
          if(_zz_2[1366]) begin
            regVec_1366 <= _zz_regVec_0_1;
          end
          if(_zz_2[1367]) begin
            regVec_1367 <= _zz_regVec_0_1;
          end
          if(_zz_2[1368]) begin
            regVec_1368 <= _zz_regVec_0_1;
          end
          if(_zz_2[1369]) begin
            regVec_1369 <= _zz_regVec_0_1;
          end
          if(_zz_2[1370]) begin
            regVec_1370 <= _zz_regVec_0_1;
          end
          if(_zz_2[1371]) begin
            regVec_1371 <= _zz_regVec_0_1;
          end
          if(_zz_2[1372]) begin
            regVec_1372 <= _zz_regVec_0_1;
          end
          if(_zz_2[1373]) begin
            regVec_1373 <= _zz_regVec_0_1;
          end
          if(_zz_2[1374]) begin
            regVec_1374 <= _zz_regVec_0_1;
          end
          if(_zz_2[1375]) begin
            regVec_1375 <= _zz_regVec_0_1;
          end
          if(_zz_2[1376]) begin
            regVec_1376 <= _zz_regVec_0_1;
          end
          if(_zz_2[1377]) begin
            regVec_1377 <= _zz_regVec_0_1;
          end
          if(_zz_2[1378]) begin
            regVec_1378 <= _zz_regVec_0_1;
          end
          if(_zz_2[1379]) begin
            regVec_1379 <= _zz_regVec_0_1;
          end
          if(_zz_2[1380]) begin
            regVec_1380 <= _zz_regVec_0_1;
          end
          if(_zz_2[1381]) begin
            regVec_1381 <= _zz_regVec_0_1;
          end
          if(_zz_2[1382]) begin
            regVec_1382 <= _zz_regVec_0_1;
          end
          if(_zz_2[1383]) begin
            regVec_1383 <= _zz_regVec_0_1;
          end
          if(_zz_2[1384]) begin
            regVec_1384 <= _zz_regVec_0_1;
          end
          if(_zz_2[1385]) begin
            regVec_1385 <= _zz_regVec_0_1;
          end
          if(_zz_2[1386]) begin
            regVec_1386 <= _zz_regVec_0_1;
          end
          if(_zz_2[1387]) begin
            regVec_1387 <= _zz_regVec_0_1;
          end
          if(_zz_2[1388]) begin
            regVec_1388 <= _zz_regVec_0_1;
          end
          if(_zz_2[1389]) begin
            regVec_1389 <= _zz_regVec_0_1;
          end
          if(_zz_2[1390]) begin
            regVec_1390 <= _zz_regVec_0_1;
          end
          if(_zz_2[1391]) begin
            regVec_1391 <= _zz_regVec_0_1;
          end
          if(_zz_2[1392]) begin
            regVec_1392 <= _zz_regVec_0_1;
          end
          if(_zz_2[1393]) begin
            regVec_1393 <= _zz_regVec_0_1;
          end
          if(_zz_2[1394]) begin
            regVec_1394 <= _zz_regVec_0_1;
          end
          if(_zz_2[1395]) begin
            regVec_1395 <= _zz_regVec_0_1;
          end
          if(_zz_2[1396]) begin
            regVec_1396 <= _zz_regVec_0_1;
          end
          if(_zz_2[1397]) begin
            regVec_1397 <= _zz_regVec_0_1;
          end
          if(_zz_2[1398]) begin
            regVec_1398 <= _zz_regVec_0_1;
          end
          if(_zz_2[1399]) begin
            regVec_1399 <= _zz_regVec_0_1;
          end
          if(_zz_2[1400]) begin
            regVec_1400 <= _zz_regVec_0_1;
          end
          if(_zz_2[1401]) begin
            regVec_1401 <= _zz_regVec_0_1;
          end
          if(_zz_2[1402]) begin
            regVec_1402 <= _zz_regVec_0_1;
          end
          if(_zz_2[1403]) begin
            regVec_1403 <= _zz_regVec_0_1;
          end
          if(_zz_2[1404]) begin
            regVec_1404 <= _zz_regVec_0_1;
          end
          if(_zz_2[1405]) begin
            regVec_1405 <= _zz_regVec_0_1;
          end
          if(_zz_2[1406]) begin
            regVec_1406 <= _zz_regVec_0_1;
          end
          if(_zz_2[1407]) begin
            regVec_1407 <= _zz_regVec_0_1;
          end
          if(_zz_2[1408]) begin
            regVec_1408 <= _zz_regVec_0_1;
          end
          if(_zz_2[1409]) begin
            regVec_1409 <= _zz_regVec_0_1;
          end
          if(_zz_2[1410]) begin
            regVec_1410 <= _zz_regVec_0_1;
          end
          if(_zz_2[1411]) begin
            regVec_1411 <= _zz_regVec_0_1;
          end
          if(_zz_2[1412]) begin
            regVec_1412 <= _zz_regVec_0_1;
          end
          if(_zz_2[1413]) begin
            regVec_1413 <= _zz_regVec_0_1;
          end
          if(_zz_2[1414]) begin
            regVec_1414 <= _zz_regVec_0_1;
          end
          if(_zz_2[1415]) begin
            regVec_1415 <= _zz_regVec_0_1;
          end
          if(_zz_2[1416]) begin
            regVec_1416 <= _zz_regVec_0_1;
          end
          if(_zz_2[1417]) begin
            regVec_1417 <= _zz_regVec_0_1;
          end
          if(_zz_2[1418]) begin
            regVec_1418 <= _zz_regVec_0_1;
          end
          if(_zz_2[1419]) begin
            regVec_1419 <= _zz_regVec_0_1;
          end
          if(_zz_2[1420]) begin
            regVec_1420 <= _zz_regVec_0_1;
          end
          if(_zz_2[1421]) begin
            regVec_1421 <= _zz_regVec_0_1;
          end
          if(_zz_2[1422]) begin
            regVec_1422 <= _zz_regVec_0_1;
          end
          if(_zz_2[1423]) begin
            regVec_1423 <= _zz_regVec_0_1;
          end
          if(_zz_2[1424]) begin
            regVec_1424 <= _zz_regVec_0_1;
          end
          if(_zz_2[1425]) begin
            regVec_1425 <= _zz_regVec_0_1;
          end
          if(_zz_2[1426]) begin
            regVec_1426 <= _zz_regVec_0_1;
          end
          if(_zz_2[1427]) begin
            regVec_1427 <= _zz_regVec_0_1;
          end
          if(_zz_2[1428]) begin
            regVec_1428 <= _zz_regVec_0_1;
          end
          if(_zz_2[1429]) begin
            regVec_1429 <= _zz_regVec_0_1;
          end
          if(_zz_2[1430]) begin
            regVec_1430 <= _zz_regVec_0_1;
          end
          if(_zz_2[1431]) begin
            regVec_1431 <= _zz_regVec_0_1;
          end
          if(_zz_2[1432]) begin
            regVec_1432 <= _zz_regVec_0_1;
          end
          if(_zz_2[1433]) begin
            regVec_1433 <= _zz_regVec_0_1;
          end
          if(_zz_2[1434]) begin
            regVec_1434 <= _zz_regVec_0_1;
          end
          if(_zz_2[1435]) begin
            regVec_1435 <= _zz_regVec_0_1;
          end
          if(_zz_2[1436]) begin
            regVec_1436 <= _zz_regVec_0_1;
          end
          if(_zz_2[1437]) begin
            regVec_1437 <= _zz_regVec_0_1;
          end
          if(_zz_2[1438]) begin
            regVec_1438 <= _zz_regVec_0_1;
          end
          if(_zz_2[1439]) begin
            regVec_1439 <= _zz_regVec_0_1;
          end
          if(_zz_2[1440]) begin
            regVec_1440 <= _zz_regVec_0_1;
          end
          if(_zz_2[1441]) begin
            regVec_1441 <= _zz_regVec_0_1;
          end
          if(_zz_2[1442]) begin
            regVec_1442 <= _zz_regVec_0_1;
          end
          if(_zz_2[1443]) begin
            regVec_1443 <= _zz_regVec_0_1;
          end
          if(_zz_2[1444]) begin
            regVec_1444 <= _zz_regVec_0_1;
          end
          if(_zz_2[1445]) begin
            regVec_1445 <= _zz_regVec_0_1;
          end
          if(_zz_2[1446]) begin
            regVec_1446 <= _zz_regVec_0_1;
          end
          if(_zz_2[1447]) begin
            regVec_1447 <= _zz_regVec_0_1;
          end
          if(_zz_2[1448]) begin
            regVec_1448 <= _zz_regVec_0_1;
          end
          if(_zz_2[1449]) begin
            regVec_1449 <= _zz_regVec_0_1;
          end
          if(_zz_2[1450]) begin
            regVec_1450 <= _zz_regVec_0_1;
          end
          if(_zz_2[1451]) begin
            regVec_1451 <= _zz_regVec_0_1;
          end
          if(_zz_2[1452]) begin
            regVec_1452 <= _zz_regVec_0_1;
          end
          if(_zz_2[1453]) begin
            regVec_1453 <= _zz_regVec_0_1;
          end
          if(_zz_2[1454]) begin
            regVec_1454 <= _zz_regVec_0_1;
          end
          if(_zz_2[1455]) begin
            regVec_1455 <= _zz_regVec_0_1;
          end
          if(_zz_2[1456]) begin
            regVec_1456 <= _zz_regVec_0_1;
          end
          if(_zz_2[1457]) begin
            regVec_1457 <= _zz_regVec_0_1;
          end
          if(_zz_2[1458]) begin
            regVec_1458 <= _zz_regVec_0_1;
          end
          if(_zz_2[1459]) begin
            regVec_1459 <= _zz_regVec_0_1;
          end
          if(_zz_2[1460]) begin
            regVec_1460 <= _zz_regVec_0_1;
          end
          if(_zz_2[1461]) begin
            regVec_1461 <= _zz_regVec_0_1;
          end
          if(_zz_2[1462]) begin
            regVec_1462 <= _zz_regVec_0_1;
          end
          if(_zz_2[1463]) begin
            regVec_1463 <= _zz_regVec_0_1;
          end
          if(_zz_2[1464]) begin
            regVec_1464 <= _zz_regVec_0_1;
          end
          if(_zz_2[1465]) begin
            regVec_1465 <= _zz_regVec_0_1;
          end
          if(_zz_2[1466]) begin
            regVec_1466 <= _zz_regVec_0_1;
          end
          if(_zz_2[1467]) begin
            regVec_1467 <= _zz_regVec_0_1;
          end
          if(_zz_2[1468]) begin
            regVec_1468 <= _zz_regVec_0_1;
          end
          if(_zz_2[1469]) begin
            regVec_1469 <= _zz_regVec_0_1;
          end
          if(_zz_2[1470]) begin
            regVec_1470 <= _zz_regVec_0_1;
          end
          if(_zz_2[1471]) begin
            regVec_1471 <= _zz_regVec_0_1;
          end
          if(_zz_2[1472]) begin
            regVec_1472 <= _zz_regVec_0_1;
          end
          if(_zz_2[1473]) begin
            regVec_1473 <= _zz_regVec_0_1;
          end
          if(_zz_2[1474]) begin
            regVec_1474 <= _zz_regVec_0_1;
          end
          if(_zz_2[1475]) begin
            regVec_1475 <= _zz_regVec_0_1;
          end
          if(_zz_2[1476]) begin
            regVec_1476 <= _zz_regVec_0_1;
          end
          if(_zz_2[1477]) begin
            regVec_1477 <= _zz_regVec_0_1;
          end
          if(_zz_2[1478]) begin
            regVec_1478 <= _zz_regVec_0_1;
          end
          if(_zz_2[1479]) begin
            regVec_1479 <= _zz_regVec_0_1;
          end
          if(_zz_2[1480]) begin
            regVec_1480 <= _zz_regVec_0_1;
          end
          if(_zz_2[1481]) begin
            regVec_1481 <= _zz_regVec_0_1;
          end
          if(_zz_2[1482]) begin
            regVec_1482 <= _zz_regVec_0_1;
          end
          if(_zz_2[1483]) begin
            regVec_1483 <= _zz_regVec_0_1;
          end
          if(_zz_2[1484]) begin
            regVec_1484 <= _zz_regVec_0_1;
          end
          if(_zz_2[1485]) begin
            regVec_1485 <= _zz_regVec_0_1;
          end
          if(_zz_2[1486]) begin
            regVec_1486 <= _zz_regVec_0_1;
          end
          if(_zz_2[1487]) begin
            regVec_1487 <= _zz_regVec_0_1;
          end
          if(_zz_2[1488]) begin
            regVec_1488 <= _zz_regVec_0_1;
          end
          if(_zz_2[1489]) begin
            regVec_1489 <= _zz_regVec_0_1;
          end
          if(_zz_2[1490]) begin
            regVec_1490 <= _zz_regVec_0_1;
          end
          if(_zz_2[1491]) begin
            regVec_1491 <= _zz_regVec_0_1;
          end
          if(_zz_2[1492]) begin
            regVec_1492 <= _zz_regVec_0_1;
          end
          if(_zz_2[1493]) begin
            regVec_1493 <= _zz_regVec_0_1;
          end
          if(_zz_2[1494]) begin
            regVec_1494 <= _zz_regVec_0_1;
          end
          if(_zz_2[1495]) begin
            regVec_1495 <= _zz_regVec_0_1;
          end
          if(_zz_2[1496]) begin
            regVec_1496 <= _zz_regVec_0_1;
          end
          if(_zz_2[1497]) begin
            regVec_1497 <= _zz_regVec_0_1;
          end
          if(_zz_2[1498]) begin
            regVec_1498 <= _zz_regVec_0_1;
          end
          if(_zz_2[1499]) begin
            regVec_1499 <= _zz_regVec_0_1;
          end
          if(_zz_2[1500]) begin
            regVec_1500 <= _zz_regVec_0_1;
          end
          if(_zz_2[1501]) begin
            regVec_1501 <= _zz_regVec_0_1;
          end
          if(_zz_2[1502]) begin
            regVec_1502 <= _zz_regVec_0_1;
          end
          if(_zz_2[1503]) begin
            regVec_1503 <= _zz_regVec_0_1;
          end
          if(_zz_2[1504]) begin
            regVec_1504 <= _zz_regVec_0_1;
          end
          if(_zz_2[1505]) begin
            regVec_1505 <= _zz_regVec_0_1;
          end
          if(_zz_2[1506]) begin
            regVec_1506 <= _zz_regVec_0_1;
          end
          if(_zz_2[1507]) begin
            regVec_1507 <= _zz_regVec_0_1;
          end
          if(_zz_2[1508]) begin
            regVec_1508 <= _zz_regVec_0_1;
          end
          if(_zz_2[1509]) begin
            regVec_1509 <= _zz_regVec_0_1;
          end
          if(_zz_2[1510]) begin
            regVec_1510 <= _zz_regVec_0_1;
          end
          if(_zz_2[1511]) begin
            regVec_1511 <= _zz_regVec_0_1;
          end
          if(_zz_2[1512]) begin
            regVec_1512 <= _zz_regVec_0_1;
          end
          if(_zz_2[1513]) begin
            regVec_1513 <= _zz_regVec_0_1;
          end
          if(_zz_2[1514]) begin
            regVec_1514 <= _zz_regVec_0_1;
          end
          if(_zz_2[1515]) begin
            regVec_1515 <= _zz_regVec_0_1;
          end
          if(_zz_2[1516]) begin
            regVec_1516 <= _zz_regVec_0_1;
          end
          if(_zz_2[1517]) begin
            regVec_1517 <= _zz_regVec_0_1;
          end
          if(_zz_2[1518]) begin
            regVec_1518 <= _zz_regVec_0_1;
          end
          if(_zz_2[1519]) begin
            regVec_1519 <= _zz_regVec_0_1;
          end
          if(_zz_2[1520]) begin
            regVec_1520 <= _zz_regVec_0_1;
          end
          if(_zz_2[1521]) begin
            regVec_1521 <= _zz_regVec_0_1;
          end
          if(_zz_2[1522]) begin
            regVec_1522 <= _zz_regVec_0_1;
          end
          if(_zz_2[1523]) begin
            regVec_1523 <= _zz_regVec_0_1;
          end
          if(_zz_2[1524]) begin
            regVec_1524 <= _zz_regVec_0_1;
          end
          if(_zz_2[1525]) begin
            regVec_1525 <= _zz_regVec_0_1;
          end
          if(_zz_2[1526]) begin
            regVec_1526 <= _zz_regVec_0_1;
          end
          if(_zz_2[1527]) begin
            regVec_1527 <= _zz_regVec_0_1;
          end
          if(_zz_2[1528]) begin
            regVec_1528 <= _zz_regVec_0_1;
          end
          if(_zz_2[1529]) begin
            regVec_1529 <= _zz_regVec_0_1;
          end
          if(_zz_2[1530]) begin
            regVec_1530 <= _zz_regVec_0_1;
          end
          if(_zz_2[1531]) begin
            regVec_1531 <= _zz_regVec_0_1;
          end
          if(_zz_2[1532]) begin
            regVec_1532 <= _zz_regVec_0_1;
          end
          if(_zz_2[1533]) begin
            regVec_1533 <= _zz_regVec_0_1;
          end
          if(_zz_2[1534]) begin
            regVec_1534 <= _zz_regVec_0_1;
          end
          if(_zz_2[1535]) begin
            regVec_1535 <= _zz_regVec_0_1;
          end
          if(_zz_2[1536]) begin
            regVec_1536 <= _zz_regVec_0_1;
          end
          if(_zz_2[1537]) begin
            regVec_1537 <= _zz_regVec_0_1;
          end
          if(_zz_2[1538]) begin
            regVec_1538 <= _zz_regVec_0_1;
          end
          if(_zz_2[1539]) begin
            regVec_1539 <= _zz_regVec_0_1;
          end
          if(_zz_2[1540]) begin
            regVec_1540 <= _zz_regVec_0_1;
          end
          if(_zz_2[1541]) begin
            regVec_1541 <= _zz_regVec_0_1;
          end
          if(_zz_2[1542]) begin
            regVec_1542 <= _zz_regVec_0_1;
          end
          if(_zz_2[1543]) begin
            regVec_1543 <= _zz_regVec_0_1;
          end
          if(_zz_2[1544]) begin
            regVec_1544 <= _zz_regVec_0_1;
          end
          if(_zz_2[1545]) begin
            regVec_1545 <= _zz_regVec_0_1;
          end
          if(_zz_2[1546]) begin
            regVec_1546 <= _zz_regVec_0_1;
          end
          if(_zz_2[1547]) begin
            regVec_1547 <= _zz_regVec_0_1;
          end
          if(_zz_2[1548]) begin
            regVec_1548 <= _zz_regVec_0_1;
          end
          if(_zz_2[1549]) begin
            regVec_1549 <= _zz_regVec_0_1;
          end
          if(_zz_2[1550]) begin
            regVec_1550 <= _zz_regVec_0_1;
          end
          if(_zz_2[1551]) begin
            regVec_1551 <= _zz_regVec_0_1;
          end
          if(_zz_2[1552]) begin
            regVec_1552 <= _zz_regVec_0_1;
          end
          if(_zz_2[1553]) begin
            regVec_1553 <= _zz_regVec_0_1;
          end
          if(_zz_2[1554]) begin
            regVec_1554 <= _zz_regVec_0_1;
          end
          if(_zz_2[1555]) begin
            regVec_1555 <= _zz_regVec_0_1;
          end
          if(_zz_2[1556]) begin
            regVec_1556 <= _zz_regVec_0_1;
          end
          if(_zz_2[1557]) begin
            regVec_1557 <= _zz_regVec_0_1;
          end
          if(_zz_2[1558]) begin
            regVec_1558 <= _zz_regVec_0_1;
          end
          if(_zz_2[1559]) begin
            regVec_1559 <= _zz_regVec_0_1;
          end
          if(_zz_2[1560]) begin
            regVec_1560 <= _zz_regVec_0_1;
          end
          if(_zz_2[1561]) begin
            regVec_1561 <= _zz_regVec_0_1;
          end
          if(_zz_2[1562]) begin
            regVec_1562 <= _zz_regVec_0_1;
          end
          if(_zz_2[1563]) begin
            regVec_1563 <= _zz_regVec_0_1;
          end
          if(_zz_2[1564]) begin
            regVec_1564 <= _zz_regVec_0_1;
          end
          if(_zz_2[1565]) begin
            regVec_1565 <= _zz_regVec_0_1;
          end
          if(_zz_2[1566]) begin
            regVec_1566 <= _zz_regVec_0_1;
          end
          if(_zz_2[1567]) begin
            regVec_1567 <= _zz_regVec_0_1;
          end
          if(_zz_2[1568]) begin
            regVec_1568 <= _zz_regVec_0_1;
          end
          if(_zz_2[1569]) begin
            regVec_1569 <= _zz_regVec_0_1;
          end
          if(_zz_2[1570]) begin
            regVec_1570 <= _zz_regVec_0_1;
          end
          if(_zz_2[1571]) begin
            regVec_1571 <= _zz_regVec_0_1;
          end
          if(_zz_2[1572]) begin
            regVec_1572 <= _zz_regVec_0_1;
          end
          if(_zz_2[1573]) begin
            regVec_1573 <= _zz_regVec_0_1;
          end
          if(_zz_2[1574]) begin
            regVec_1574 <= _zz_regVec_0_1;
          end
          if(_zz_2[1575]) begin
            regVec_1575 <= _zz_regVec_0_1;
          end
          if(_zz_2[1576]) begin
            regVec_1576 <= _zz_regVec_0_1;
          end
          if(_zz_2[1577]) begin
            regVec_1577 <= _zz_regVec_0_1;
          end
          if(_zz_2[1578]) begin
            regVec_1578 <= _zz_regVec_0_1;
          end
          if(_zz_2[1579]) begin
            regVec_1579 <= _zz_regVec_0_1;
          end
          if(_zz_2[1580]) begin
            regVec_1580 <= _zz_regVec_0_1;
          end
          if(_zz_2[1581]) begin
            regVec_1581 <= _zz_regVec_0_1;
          end
          if(_zz_2[1582]) begin
            regVec_1582 <= _zz_regVec_0_1;
          end
          if(_zz_2[1583]) begin
            regVec_1583 <= _zz_regVec_0_1;
          end
          if(_zz_2[1584]) begin
            regVec_1584 <= _zz_regVec_0_1;
          end
          if(_zz_2[1585]) begin
            regVec_1585 <= _zz_regVec_0_1;
          end
          if(_zz_2[1586]) begin
            regVec_1586 <= _zz_regVec_0_1;
          end
          if(_zz_2[1587]) begin
            regVec_1587 <= _zz_regVec_0_1;
          end
          if(_zz_2[1588]) begin
            regVec_1588 <= _zz_regVec_0_1;
          end
          if(_zz_2[1589]) begin
            regVec_1589 <= _zz_regVec_0_1;
          end
          if(_zz_2[1590]) begin
            regVec_1590 <= _zz_regVec_0_1;
          end
          if(_zz_2[1591]) begin
            regVec_1591 <= _zz_regVec_0_1;
          end
          if(_zz_2[1592]) begin
            regVec_1592 <= _zz_regVec_0_1;
          end
          if(_zz_2[1593]) begin
            regVec_1593 <= _zz_regVec_0_1;
          end
          if(_zz_2[1594]) begin
            regVec_1594 <= _zz_regVec_0_1;
          end
          if(_zz_2[1595]) begin
            regVec_1595 <= _zz_regVec_0_1;
          end
          if(_zz_2[1596]) begin
            regVec_1596 <= _zz_regVec_0_1;
          end
          if(_zz_2[1597]) begin
            regVec_1597 <= _zz_regVec_0_1;
          end
          if(_zz_2[1598]) begin
            regVec_1598 <= _zz_regVec_0_1;
          end
          if(_zz_2[1599]) begin
            regVec_1599 <= _zz_regVec_0_1;
          end
          if(_zz_2[1600]) begin
            regVec_1600 <= _zz_regVec_0_1;
          end
          if(_zz_2[1601]) begin
            regVec_1601 <= _zz_regVec_0_1;
          end
          if(_zz_2[1602]) begin
            regVec_1602 <= _zz_regVec_0_1;
          end
          if(_zz_2[1603]) begin
            regVec_1603 <= _zz_regVec_0_1;
          end
          if(_zz_2[1604]) begin
            regVec_1604 <= _zz_regVec_0_1;
          end
          if(_zz_2[1605]) begin
            regVec_1605 <= _zz_regVec_0_1;
          end
          if(_zz_2[1606]) begin
            regVec_1606 <= _zz_regVec_0_1;
          end
          if(_zz_2[1607]) begin
            regVec_1607 <= _zz_regVec_0_1;
          end
          if(_zz_2[1608]) begin
            regVec_1608 <= _zz_regVec_0_1;
          end
          if(_zz_2[1609]) begin
            regVec_1609 <= _zz_regVec_0_1;
          end
          if(_zz_2[1610]) begin
            regVec_1610 <= _zz_regVec_0_1;
          end
          if(_zz_2[1611]) begin
            regVec_1611 <= _zz_regVec_0_1;
          end
          if(_zz_2[1612]) begin
            regVec_1612 <= _zz_regVec_0_1;
          end
          if(_zz_2[1613]) begin
            regVec_1613 <= _zz_regVec_0_1;
          end
          if(_zz_2[1614]) begin
            regVec_1614 <= _zz_regVec_0_1;
          end
          if(_zz_2[1615]) begin
            regVec_1615 <= _zz_regVec_0_1;
          end
          if(_zz_2[1616]) begin
            regVec_1616 <= _zz_regVec_0_1;
          end
          if(_zz_2[1617]) begin
            regVec_1617 <= _zz_regVec_0_1;
          end
          if(_zz_2[1618]) begin
            regVec_1618 <= _zz_regVec_0_1;
          end
          if(_zz_2[1619]) begin
            regVec_1619 <= _zz_regVec_0_1;
          end
          if(_zz_2[1620]) begin
            regVec_1620 <= _zz_regVec_0_1;
          end
          if(_zz_2[1621]) begin
            regVec_1621 <= _zz_regVec_0_1;
          end
          if(_zz_2[1622]) begin
            regVec_1622 <= _zz_regVec_0_1;
          end
          if(_zz_2[1623]) begin
            regVec_1623 <= _zz_regVec_0_1;
          end
          if(_zz_2[1624]) begin
            regVec_1624 <= _zz_regVec_0_1;
          end
          if(_zz_2[1625]) begin
            regVec_1625 <= _zz_regVec_0_1;
          end
          if(_zz_2[1626]) begin
            regVec_1626 <= _zz_regVec_0_1;
          end
          if(_zz_2[1627]) begin
            regVec_1627 <= _zz_regVec_0_1;
          end
          if(_zz_2[1628]) begin
            regVec_1628 <= _zz_regVec_0_1;
          end
          if(_zz_2[1629]) begin
            regVec_1629 <= _zz_regVec_0_1;
          end
          if(_zz_2[1630]) begin
            regVec_1630 <= _zz_regVec_0_1;
          end
          if(_zz_2[1631]) begin
            regVec_1631 <= _zz_regVec_0_1;
          end
          if(_zz_2[1632]) begin
            regVec_1632 <= _zz_regVec_0_1;
          end
          if(_zz_2[1633]) begin
            regVec_1633 <= _zz_regVec_0_1;
          end
          if(_zz_2[1634]) begin
            regVec_1634 <= _zz_regVec_0_1;
          end
          if(_zz_2[1635]) begin
            regVec_1635 <= _zz_regVec_0_1;
          end
          if(_zz_2[1636]) begin
            regVec_1636 <= _zz_regVec_0_1;
          end
          if(_zz_2[1637]) begin
            regVec_1637 <= _zz_regVec_0_1;
          end
          if(_zz_2[1638]) begin
            regVec_1638 <= _zz_regVec_0_1;
          end
          if(_zz_2[1639]) begin
            regVec_1639 <= _zz_regVec_0_1;
          end
          if(_zz_2[1640]) begin
            regVec_1640 <= _zz_regVec_0_1;
          end
          if(_zz_2[1641]) begin
            regVec_1641 <= _zz_regVec_0_1;
          end
          if(_zz_2[1642]) begin
            regVec_1642 <= _zz_regVec_0_1;
          end
          if(_zz_2[1643]) begin
            regVec_1643 <= _zz_regVec_0_1;
          end
          if(_zz_2[1644]) begin
            regVec_1644 <= _zz_regVec_0_1;
          end
          if(_zz_2[1645]) begin
            regVec_1645 <= _zz_regVec_0_1;
          end
          if(_zz_2[1646]) begin
            regVec_1646 <= _zz_regVec_0_1;
          end
          if(_zz_2[1647]) begin
            regVec_1647 <= _zz_regVec_0_1;
          end
          if(_zz_2[1648]) begin
            regVec_1648 <= _zz_regVec_0_1;
          end
          if(_zz_2[1649]) begin
            regVec_1649 <= _zz_regVec_0_1;
          end
          if(_zz_2[1650]) begin
            regVec_1650 <= _zz_regVec_0_1;
          end
          if(_zz_2[1651]) begin
            regVec_1651 <= _zz_regVec_0_1;
          end
          if(_zz_2[1652]) begin
            regVec_1652 <= _zz_regVec_0_1;
          end
          if(_zz_2[1653]) begin
            regVec_1653 <= _zz_regVec_0_1;
          end
          if(_zz_2[1654]) begin
            regVec_1654 <= _zz_regVec_0_1;
          end
          if(_zz_2[1655]) begin
            regVec_1655 <= _zz_regVec_0_1;
          end
          if(_zz_2[1656]) begin
            regVec_1656 <= _zz_regVec_0_1;
          end
          if(_zz_2[1657]) begin
            regVec_1657 <= _zz_regVec_0_1;
          end
          if(_zz_2[1658]) begin
            regVec_1658 <= _zz_regVec_0_1;
          end
          if(_zz_2[1659]) begin
            regVec_1659 <= _zz_regVec_0_1;
          end
          if(_zz_2[1660]) begin
            regVec_1660 <= _zz_regVec_0_1;
          end
          if(_zz_2[1661]) begin
            regVec_1661 <= _zz_regVec_0_1;
          end
          if(_zz_2[1662]) begin
            regVec_1662 <= _zz_regVec_0_1;
          end
          if(_zz_2[1663]) begin
            regVec_1663 <= _zz_regVec_0_1;
          end
          if(_zz_2[1664]) begin
            regVec_1664 <= _zz_regVec_0_1;
          end
          if(_zz_2[1665]) begin
            regVec_1665 <= _zz_regVec_0_1;
          end
          if(_zz_2[1666]) begin
            regVec_1666 <= _zz_regVec_0_1;
          end
          if(_zz_2[1667]) begin
            regVec_1667 <= _zz_regVec_0_1;
          end
          if(_zz_2[1668]) begin
            regVec_1668 <= _zz_regVec_0_1;
          end
          if(_zz_2[1669]) begin
            regVec_1669 <= _zz_regVec_0_1;
          end
          if(_zz_2[1670]) begin
            regVec_1670 <= _zz_regVec_0_1;
          end
          if(_zz_2[1671]) begin
            regVec_1671 <= _zz_regVec_0_1;
          end
          if(_zz_2[1672]) begin
            regVec_1672 <= _zz_regVec_0_1;
          end
          if(_zz_2[1673]) begin
            regVec_1673 <= _zz_regVec_0_1;
          end
          if(_zz_2[1674]) begin
            regVec_1674 <= _zz_regVec_0_1;
          end
          if(_zz_2[1675]) begin
            regVec_1675 <= _zz_regVec_0_1;
          end
          if(_zz_2[1676]) begin
            regVec_1676 <= _zz_regVec_0_1;
          end
          if(_zz_2[1677]) begin
            regVec_1677 <= _zz_regVec_0_1;
          end
          if(_zz_2[1678]) begin
            regVec_1678 <= _zz_regVec_0_1;
          end
          if(_zz_2[1679]) begin
            regVec_1679 <= _zz_regVec_0_1;
          end
          if(_zz_2[1680]) begin
            regVec_1680 <= _zz_regVec_0_1;
          end
          if(_zz_2[1681]) begin
            regVec_1681 <= _zz_regVec_0_1;
          end
          if(_zz_2[1682]) begin
            regVec_1682 <= _zz_regVec_0_1;
          end
          if(_zz_2[1683]) begin
            regVec_1683 <= _zz_regVec_0_1;
          end
          if(_zz_2[1684]) begin
            regVec_1684 <= _zz_regVec_0_1;
          end
          if(_zz_2[1685]) begin
            regVec_1685 <= _zz_regVec_0_1;
          end
          if(_zz_2[1686]) begin
            regVec_1686 <= _zz_regVec_0_1;
          end
          if(_zz_2[1687]) begin
            regVec_1687 <= _zz_regVec_0_1;
          end
          if(_zz_2[1688]) begin
            regVec_1688 <= _zz_regVec_0_1;
          end
          if(_zz_2[1689]) begin
            regVec_1689 <= _zz_regVec_0_1;
          end
          if(_zz_2[1690]) begin
            regVec_1690 <= _zz_regVec_0_1;
          end
          if(_zz_2[1691]) begin
            regVec_1691 <= _zz_regVec_0_1;
          end
          if(_zz_2[1692]) begin
            regVec_1692 <= _zz_regVec_0_1;
          end
          if(_zz_2[1693]) begin
            regVec_1693 <= _zz_regVec_0_1;
          end
          if(_zz_2[1694]) begin
            regVec_1694 <= _zz_regVec_0_1;
          end
          if(_zz_2[1695]) begin
            regVec_1695 <= _zz_regVec_0_1;
          end
          if(_zz_2[1696]) begin
            regVec_1696 <= _zz_regVec_0_1;
          end
          if(_zz_2[1697]) begin
            regVec_1697 <= _zz_regVec_0_1;
          end
          if(_zz_2[1698]) begin
            regVec_1698 <= _zz_regVec_0_1;
          end
          if(_zz_2[1699]) begin
            regVec_1699 <= _zz_regVec_0_1;
          end
          if(_zz_2[1700]) begin
            regVec_1700 <= _zz_regVec_0_1;
          end
          if(_zz_2[1701]) begin
            regVec_1701 <= _zz_regVec_0_1;
          end
          if(_zz_2[1702]) begin
            regVec_1702 <= _zz_regVec_0_1;
          end
          if(_zz_2[1703]) begin
            regVec_1703 <= _zz_regVec_0_1;
          end
          if(_zz_2[1704]) begin
            regVec_1704 <= _zz_regVec_0_1;
          end
          if(_zz_2[1705]) begin
            regVec_1705 <= _zz_regVec_0_1;
          end
          if(_zz_2[1706]) begin
            regVec_1706 <= _zz_regVec_0_1;
          end
          if(_zz_2[1707]) begin
            regVec_1707 <= _zz_regVec_0_1;
          end
          if(_zz_2[1708]) begin
            regVec_1708 <= _zz_regVec_0_1;
          end
          if(_zz_2[1709]) begin
            regVec_1709 <= _zz_regVec_0_1;
          end
          if(_zz_2[1710]) begin
            regVec_1710 <= _zz_regVec_0_1;
          end
          if(_zz_2[1711]) begin
            regVec_1711 <= _zz_regVec_0_1;
          end
          if(_zz_2[1712]) begin
            regVec_1712 <= _zz_regVec_0_1;
          end
          if(_zz_2[1713]) begin
            regVec_1713 <= _zz_regVec_0_1;
          end
          if(_zz_2[1714]) begin
            regVec_1714 <= _zz_regVec_0_1;
          end
          if(_zz_2[1715]) begin
            regVec_1715 <= _zz_regVec_0_1;
          end
          if(_zz_2[1716]) begin
            regVec_1716 <= _zz_regVec_0_1;
          end
          if(_zz_2[1717]) begin
            regVec_1717 <= _zz_regVec_0_1;
          end
          if(_zz_2[1718]) begin
            regVec_1718 <= _zz_regVec_0_1;
          end
          if(_zz_2[1719]) begin
            regVec_1719 <= _zz_regVec_0_1;
          end
          if(_zz_2[1720]) begin
            regVec_1720 <= _zz_regVec_0_1;
          end
          if(_zz_2[1721]) begin
            regVec_1721 <= _zz_regVec_0_1;
          end
          if(_zz_2[1722]) begin
            regVec_1722 <= _zz_regVec_0_1;
          end
          if(_zz_2[1723]) begin
            regVec_1723 <= _zz_regVec_0_1;
          end
          if(_zz_2[1724]) begin
            regVec_1724 <= _zz_regVec_0_1;
          end
          if(_zz_2[1725]) begin
            regVec_1725 <= _zz_regVec_0_1;
          end
          if(_zz_2[1726]) begin
            regVec_1726 <= _zz_regVec_0_1;
          end
          if(_zz_2[1727]) begin
            regVec_1727 <= _zz_regVec_0_1;
          end
          if(_zz_2[1728]) begin
            regVec_1728 <= _zz_regVec_0_1;
          end
          if(_zz_2[1729]) begin
            regVec_1729 <= _zz_regVec_0_1;
          end
          if(_zz_2[1730]) begin
            regVec_1730 <= _zz_regVec_0_1;
          end
          if(_zz_2[1731]) begin
            regVec_1731 <= _zz_regVec_0_1;
          end
          if(_zz_2[1732]) begin
            regVec_1732 <= _zz_regVec_0_1;
          end
          if(_zz_2[1733]) begin
            regVec_1733 <= _zz_regVec_0_1;
          end
          if(_zz_2[1734]) begin
            regVec_1734 <= _zz_regVec_0_1;
          end
          if(_zz_2[1735]) begin
            regVec_1735 <= _zz_regVec_0_1;
          end
          if(_zz_2[1736]) begin
            regVec_1736 <= _zz_regVec_0_1;
          end
          if(_zz_2[1737]) begin
            regVec_1737 <= _zz_regVec_0_1;
          end
          if(_zz_2[1738]) begin
            regVec_1738 <= _zz_regVec_0_1;
          end
          if(_zz_2[1739]) begin
            regVec_1739 <= _zz_regVec_0_1;
          end
          if(_zz_2[1740]) begin
            regVec_1740 <= _zz_regVec_0_1;
          end
          if(_zz_2[1741]) begin
            regVec_1741 <= _zz_regVec_0_1;
          end
          if(_zz_2[1742]) begin
            regVec_1742 <= _zz_regVec_0_1;
          end
          if(_zz_2[1743]) begin
            regVec_1743 <= _zz_regVec_0_1;
          end
          if(_zz_2[1744]) begin
            regVec_1744 <= _zz_regVec_0_1;
          end
          if(_zz_2[1745]) begin
            regVec_1745 <= _zz_regVec_0_1;
          end
          if(_zz_2[1746]) begin
            regVec_1746 <= _zz_regVec_0_1;
          end
          if(_zz_2[1747]) begin
            regVec_1747 <= _zz_regVec_0_1;
          end
          if(_zz_2[1748]) begin
            regVec_1748 <= _zz_regVec_0_1;
          end
          if(_zz_2[1749]) begin
            regVec_1749 <= _zz_regVec_0_1;
          end
          if(_zz_2[1750]) begin
            regVec_1750 <= _zz_regVec_0_1;
          end
          if(_zz_2[1751]) begin
            regVec_1751 <= _zz_regVec_0_1;
          end
          if(_zz_2[1752]) begin
            regVec_1752 <= _zz_regVec_0_1;
          end
          if(_zz_2[1753]) begin
            regVec_1753 <= _zz_regVec_0_1;
          end
          if(_zz_2[1754]) begin
            regVec_1754 <= _zz_regVec_0_1;
          end
          if(_zz_2[1755]) begin
            regVec_1755 <= _zz_regVec_0_1;
          end
          if(_zz_2[1756]) begin
            regVec_1756 <= _zz_regVec_0_1;
          end
          if(_zz_2[1757]) begin
            regVec_1757 <= _zz_regVec_0_1;
          end
          if(_zz_2[1758]) begin
            regVec_1758 <= _zz_regVec_0_1;
          end
          if(_zz_2[1759]) begin
            regVec_1759 <= _zz_regVec_0_1;
          end
          if(_zz_2[1760]) begin
            regVec_1760 <= _zz_regVec_0_1;
          end
          if(_zz_2[1761]) begin
            regVec_1761 <= _zz_regVec_0_1;
          end
          if(_zz_2[1762]) begin
            regVec_1762 <= _zz_regVec_0_1;
          end
          if(_zz_2[1763]) begin
            regVec_1763 <= _zz_regVec_0_1;
          end
          if(_zz_2[1764]) begin
            regVec_1764 <= _zz_regVec_0_1;
          end
          if(_zz_2[1765]) begin
            regVec_1765 <= _zz_regVec_0_1;
          end
          if(_zz_2[1766]) begin
            regVec_1766 <= _zz_regVec_0_1;
          end
          if(_zz_2[1767]) begin
            regVec_1767 <= _zz_regVec_0_1;
          end
          if(_zz_2[1768]) begin
            regVec_1768 <= _zz_regVec_0_1;
          end
          if(_zz_2[1769]) begin
            regVec_1769 <= _zz_regVec_0_1;
          end
          if(_zz_2[1770]) begin
            regVec_1770 <= _zz_regVec_0_1;
          end
          if(_zz_2[1771]) begin
            regVec_1771 <= _zz_regVec_0_1;
          end
          if(_zz_2[1772]) begin
            regVec_1772 <= _zz_regVec_0_1;
          end
          if(_zz_2[1773]) begin
            regVec_1773 <= _zz_regVec_0_1;
          end
          if(_zz_2[1774]) begin
            regVec_1774 <= _zz_regVec_0_1;
          end
          if(_zz_2[1775]) begin
            regVec_1775 <= _zz_regVec_0_1;
          end
          if(_zz_2[1776]) begin
            regVec_1776 <= _zz_regVec_0_1;
          end
          if(_zz_2[1777]) begin
            regVec_1777 <= _zz_regVec_0_1;
          end
          if(_zz_2[1778]) begin
            regVec_1778 <= _zz_regVec_0_1;
          end
          if(_zz_2[1779]) begin
            regVec_1779 <= _zz_regVec_0_1;
          end
          if(_zz_2[1780]) begin
            regVec_1780 <= _zz_regVec_0_1;
          end
          if(_zz_2[1781]) begin
            regVec_1781 <= _zz_regVec_0_1;
          end
          if(_zz_2[1782]) begin
            regVec_1782 <= _zz_regVec_0_1;
          end
          if(_zz_2[1783]) begin
            regVec_1783 <= _zz_regVec_0_1;
          end
          if(_zz_2[1784]) begin
            regVec_1784 <= _zz_regVec_0_1;
          end
          if(_zz_2[1785]) begin
            regVec_1785 <= _zz_regVec_0_1;
          end
          if(_zz_2[1786]) begin
            regVec_1786 <= _zz_regVec_0_1;
          end
          if(_zz_2[1787]) begin
            regVec_1787 <= _zz_regVec_0_1;
          end
          if(_zz_2[1788]) begin
            regVec_1788 <= _zz_regVec_0_1;
          end
          if(_zz_2[1789]) begin
            regVec_1789 <= _zz_regVec_0_1;
          end
          if(_zz_2[1790]) begin
            regVec_1790 <= _zz_regVec_0_1;
          end
          if(_zz_2[1791]) begin
            regVec_1791 <= _zz_regVec_0_1;
          end
          if(_zz_2[1792]) begin
            regVec_1792 <= _zz_regVec_0_1;
          end
          if(_zz_2[1793]) begin
            regVec_1793 <= _zz_regVec_0_1;
          end
          if(_zz_2[1794]) begin
            regVec_1794 <= _zz_regVec_0_1;
          end
          if(_zz_2[1795]) begin
            regVec_1795 <= _zz_regVec_0_1;
          end
          if(_zz_2[1796]) begin
            regVec_1796 <= _zz_regVec_0_1;
          end
          if(_zz_2[1797]) begin
            regVec_1797 <= _zz_regVec_0_1;
          end
          if(_zz_2[1798]) begin
            regVec_1798 <= _zz_regVec_0_1;
          end
          if(_zz_2[1799]) begin
            regVec_1799 <= _zz_regVec_0_1;
          end
          if(_zz_2[1800]) begin
            regVec_1800 <= _zz_regVec_0_1;
          end
          if(_zz_2[1801]) begin
            regVec_1801 <= _zz_regVec_0_1;
          end
          if(_zz_2[1802]) begin
            regVec_1802 <= _zz_regVec_0_1;
          end
          if(_zz_2[1803]) begin
            regVec_1803 <= _zz_regVec_0_1;
          end
          if(_zz_2[1804]) begin
            regVec_1804 <= _zz_regVec_0_1;
          end
          if(_zz_2[1805]) begin
            regVec_1805 <= _zz_regVec_0_1;
          end
          if(_zz_2[1806]) begin
            regVec_1806 <= _zz_regVec_0_1;
          end
          if(_zz_2[1807]) begin
            regVec_1807 <= _zz_regVec_0_1;
          end
          if(_zz_2[1808]) begin
            regVec_1808 <= _zz_regVec_0_1;
          end
          if(_zz_2[1809]) begin
            regVec_1809 <= _zz_regVec_0_1;
          end
          if(_zz_2[1810]) begin
            regVec_1810 <= _zz_regVec_0_1;
          end
          if(_zz_2[1811]) begin
            regVec_1811 <= _zz_regVec_0_1;
          end
          if(_zz_2[1812]) begin
            regVec_1812 <= _zz_regVec_0_1;
          end
          if(_zz_2[1813]) begin
            regVec_1813 <= _zz_regVec_0_1;
          end
          if(_zz_2[1814]) begin
            regVec_1814 <= _zz_regVec_0_1;
          end
          if(_zz_2[1815]) begin
            regVec_1815 <= _zz_regVec_0_1;
          end
          if(_zz_2[1816]) begin
            regVec_1816 <= _zz_regVec_0_1;
          end
          if(_zz_2[1817]) begin
            regVec_1817 <= _zz_regVec_0_1;
          end
          if(_zz_2[1818]) begin
            regVec_1818 <= _zz_regVec_0_1;
          end
          if(_zz_2[1819]) begin
            regVec_1819 <= _zz_regVec_0_1;
          end
          if(_zz_2[1820]) begin
            regVec_1820 <= _zz_regVec_0_1;
          end
          if(_zz_2[1821]) begin
            regVec_1821 <= _zz_regVec_0_1;
          end
          if(_zz_2[1822]) begin
            regVec_1822 <= _zz_regVec_0_1;
          end
          if(_zz_2[1823]) begin
            regVec_1823 <= _zz_regVec_0_1;
          end
          if(_zz_2[1824]) begin
            regVec_1824 <= _zz_regVec_0_1;
          end
          if(_zz_2[1825]) begin
            regVec_1825 <= _zz_regVec_0_1;
          end
          if(_zz_2[1826]) begin
            regVec_1826 <= _zz_regVec_0_1;
          end
          if(_zz_2[1827]) begin
            regVec_1827 <= _zz_regVec_0_1;
          end
          if(_zz_2[1828]) begin
            regVec_1828 <= _zz_regVec_0_1;
          end
          if(_zz_2[1829]) begin
            regVec_1829 <= _zz_regVec_0_1;
          end
          if(_zz_2[1830]) begin
            regVec_1830 <= _zz_regVec_0_1;
          end
          if(_zz_2[1831]) begin
            regVec_1831 <= _zz_regVec_0_1;
          end
          if(_zz_2[1832]) begin
            regVec_1832 <= _zz_regVec_0_1;
          end
          if(_zz_2[1833]) begin
            regVec_1833 <= _zz_regVec_0_1;
          end
          if(_zz_2[1834]) begin
            regVec_1834 <= _zz_regVec_0_1;
          end
          if(_zz_2[1835]) begin
            regVec_1835 <= _zz_regVec_0_1;
          end
          if(_zz_2[1836]) begin
            regVec_1836 <= _zz_regVec_0_1;
          end
          if(_zz_2[1837]) begin
            regVec_1837 <= _zz_regVec_0_1;
          end
          if(_zz_2[1838]) begin
            regVec_1838 <= _zz_regVec_0_1;
          end
          if(_zz_2[1839]) begin
            regVec_1839 <= _zz_regVec_0_1;
          end
          if(_zz_2[1840]) begin
            regVec_1840 <= _zz_regVec_0_1;
          end
          if(_zz_2[1841]) begin
            regVec_1841 <= _zz_regVec_0_1;
          end
          if(_zz_2[1842]) begin
            regVec_1842 <= _zz_regVec_0_1;
          end
          if(_zz_2[1843]) begin
            regVec_1843 <= _zz_regVec_0_1;
          end
          if(_zz_2[1844]) begin
            regVec_1844 <= _zz_regVec_0_1;
          end
          if(_zz_2[1845]) begin
            regVec_1845 <= _zz_regVec_0_1;
          end
          if(_zz_2[1846]) begin
            regVec_1846 <= _zz_regVec_0_1;
          end
          if(_zz_2[1847]) begin
            regVec_1847 <= _zz_regVec_0_1;
          end
          if(_zz_2[1848]) begin
            regVec_1848 <= _zz_regVec_0_1;
          end
          if(_zz_2[1849]) begin
            regVec_1849 <= _zz_regVec_0_1;
          end
          if(_zz_2[1850]) begin
            regVec_1850 <= _zz_regVec_0_1;
          end
          if(_zz_2[1851]) begin
            regVec_1851 <= _zz_regVec_0_1;
          end
          if(_zz_2[1852]) begin
            regVec_1852 <= _zz_regVec_0_1;
          end
          if(_zz_2[1853]) begin
            regVec_1853 <= _zz_regVec_0_1;
          end
          if(_zz_2[1854]) begin
            regVec_1854 <= _zz_regVec_0_1;
          end
          if(_zz_2[1855]) begin
            regVec_1855 <= _zz_regVec_0_1;
          end
          if(_zz_2[1856]) begin
            regVec_1856 <= _zz_regVec_0_1;
          end
          if(_zz_2[1857]) begin
            regVec_1857 <= _zz_regVec_0_1;
          end
          if(_zz_2[1858]) begin
            regVec_1858 <= _zz_regVec_0_1;
          end
          if(_zz_2[1859]) begin
            regVec_1859 <= _zz_regVec_0_1;
          end
          if(_zz_2[1860]) begin
            regVec_1860 <= _zz_regVec_0_1;
          end
          if(_zz_2[1861]) begin
            regVec_1861 <= _zz_regVec_0_1;
          end
          if(_zz_2[1862]) begin
            regVec_1862 <= _zz_regVec_0_1;
          end
          if(_zz_2[1863]) begin
            regVec_1863 <= _zz_regVec_0_1;
          end
          if(_zz_2[1864]) begin
            regVec_1864 <= _zz_regVec_0_1;
          end
          if(_zz_2[1865]) begin
            regVec_1865 <= _zz_regVec_0_1;
          end
          if(_zz_2[1866]) begin
            regVec_1866 <= _zz_regVec_0_1;
          end
          if(_zz_2[1867]) begin
            regVec_1867 <= _zz_regVec_0_1;
          end
          if(_zz_2[1868]) begin
            regVec_1868 <= _zz_regVec_0_1;
          end
          if(_zz_2[1869]) begin
            regVec_1869 <= _zz_regVec_0_1;
          end
          if(_zz_2[1870]) begin
            regVec_1870 <= _zz_regVec_0_1;
          end
          if(_zz_2[1871]) begin
            regVec_1871 <= _zz_regVec_0_1;
          end
          if(_zz_2[1872]) begin
            regVec_1872 <= _zz_regVec_0_1;
          end
          if(_zz_2[1873]) begin
            regVec_1873 <= _zz_regVec_0_1;
          end
          if(_zz_2[1874]) begin
            regVec_1874 <= _zz_regVec_0_1;
          end
          if(_zz_2[1875]) begin
            regVec_1875 <= _zz_regVec_0_1;
          end
          if(_zz_2[1876]) begin
            regVec_1876 <= _zz_regVec_0_1;
          end
          if(_zz_2[1877]) begin
            regVec_1877 <= _zz_regVec_0_1;
          end
          if(_zz_2[1878]) begin
            regVec_1878 <= _zz_regVec_0_1;
          end
          if(_zz_2[1879]) begin
            regVec_1879 <= _zz_regVec_0_1;
          end
          if(_zz_2[1880]) begin
            regVec_1880 <= _zz_regVec_0_1;
          end
          if(_zz_2[1881]) begin
            regVec_1881 <= _zz_regVec_0_1;
          end
          if(_zz_2[1882]) begin
            regVec_1882 <= _zz_regVec_0_1;
          end
          if(_zz_2[1883]) begin
            regVec_1883 <= _zz_regVec_0_1;
          end
          if(_zz_2[1884]) begin
            regVec_1884 <= _zz_regVec_0_1;
          end
          if(_zz_2[1885]) begin
            regVec_1885 <= _zz_regVec_0_1;
          end
          if(_zz_2[1886]) begin
            regVec_1886 <= _zz_regVec_0_1;
          end
          if(_zz_2[1887]) begin
            regVec_1887 <= _zz_regVec_0_1;
          end
          if(_zz_2[1888]) begin
            regVec_1888 <= _zz_regVec_0_1;
          end
          if(_zz_2[1889]) begin
            regVec_1889 <= _zz_regVec_0_1;
          end
          if(_zz_2[1890]) begin
            regVec_1890 <= _zz_regVec_0_1;
          end
          if(_zz_2[1891]) begin
            regVec_1891 <= _zz_regVec_0_1;
          end
          if(_zz_2[1892]) begin
            regVec_1892 <= _zz_regVec_0_1;
          end
          if(_zz_2[1893]) begin
            regVec_1893 <= _zz_regVec_0_1;
          end
          if(_zz_2[1894]) begin
            regVec_1894 <= _zz_regVec_0_1;
          end
          if(_zz_2[1895]) begin
            regVec_1895 <= _zz_regVec_0_1;
          end
          if(_zz_2[1896]) begin
            regVec_1896 <= _zz_regVec_0_1;
          end
          if(_zz_2[1897]) begin
            regVec_1897 <= _zz_regVec_0_1;
          end
          if(_zz_2[1898]) begin
            regVec_1898 <= _zz_regVec_0_1;
          end
          if(_zz_2[1899]) begin
            regVec_1899 <= _zz_regVec_0_1;
          end
          if(_zz_2[1900]) begin
            regVec_1900 <= _zz_regVec_0_1;
          end
          if(_zz_2[1901]) begin
            regVec_1901 <= _zz_regVec_0_1;
          end
          if(_zz_2[1902]) begin
            regVec_1902 <= _zz_regVec_0_1;
          end
          if(_zz_2[1903]) begin
            regVec_1903 <= _zz_regVec_0_1;
          end
          if(_zz_2[1904]) begin
            regVec_1904 <= _zz_regVec_0_1;
          end
          if(_zz_2[1905]) begin
            regVec_1905 <= _zz_regVec_0_1;
          end
          if(_zz_2[1906]) begin
            regVec_1906 <= _zz_regVec_0_1;
          end
          if(_zz_2[1907]) begin
            regVec_1907 <= _zz_regVec_0_1;
          end
          if(_zz_2[1908]) begin
            regVec_1908 <= _zz_regVec_0_1;
          end
          if(_zz_2[1909]) begin
            regVec_1909 <= _zz_regVec_0_1;
          end
          if(_zz_2[1910]) begin
            regVec_1910 <= _zz_regVec_0_1;
          end
          if(_zz_2[1911]) begin
            regVec_1911 <= _zz_regVec_0_1;
          end
          if(_zz_2[1912]) begin
            regVec_1912 <= _zz_regVec_0_1;
          end
          if(_zz_2[1913]) begin
            regVec_1913 <= _zz_regVec_0_1;
          end
          if(_zz_2[1914]) begin
            regVec_1914 <= _zz_regVec_0_1;
          end
          if(_zz_2[1915]) begin
            regVec_1915 <= _zz_regVec_0_1;
          end
          if(_zz_2[1916]) begin
            regVec_1916 <= _zz_regVec_0_1;
          end
          if(_zz_2[1917]) begin
            regVec_1917 <= _zz_regVec_0_1;
          end
          if(_zz_2[1918]) begin
            regVec_1918 <= _zz_regVec_0_1;
          end
          if(_zz_2[1919]) begin
            regVec_1919 <= _zz_regVec_0_1;
          end
          if(_zz_2[1920]) begin
            regVec_1920 <= _zz_regVec_0_1;
          end
          if(_zz_2[1921]) begin
            regVec_1921 <= _zz_regVec_0_1;
          end
          if(_zz_2[1922]) begin
            regVec_1922 <= _zz_regVec_0_1;
          end
          if(_zz_2[1923]) begin
            regVec_1923 <= _zz_regVec_0_1;
          end
          if(_zz_2[1924]) begin
            regVec_1924 <= _zz_regVec_0_1;
          end
          if(_zz_2[1925]) begin
            regVec_1925 <= _zz_regVec_0_1;
          end
          if(_zz_2[1926]) begin
            regVec_1926 <= _zz_regVec_0_1;
          end
          if(_zz_2[1927]) begin
            regVec_1927 <= _zz_regVec_0_1;
          end
          if(_zz_2[1928]) begin
            regVec_1928 <= _zz_regVec_0_1;
          end
          if(_zz_2[1929]) begin
            regVec_1929 <= _zz_regVec_0_1;
          end
          if(_zz_2[1930]) begin
            regVec_1930 <= _zz_regVec_0_1;
          end
          if(_zz_2[1931]) begin
            regVec_1931 <= _zz_regVec_0_1;
          end
          if(_zz_2[1932]) begin
            regVec_1932 <= _zz_regVec_0_1;
          end
          if(_zz_2[1933]) begin
            regVec_1933 <= _zz_regVec_0_1;
          end
          if(_zz_2[1934]) begin
            regVec_1934 <= _zz_regVec_0_1;
          end
          if(_zz_2[1935]) begin
            regVec_1935 <= _zz_regVec_0_1;
          end
          if(_zz_2[1936]) begin
            regVec_1936 <= _zz_regVec_0_1;
          end
          if(_zz_2[1937]) begin
            regVec_1937 <= _zz_regVec_0_1;
          end
          if(_zz_2[1938]) begin
            regVec_1938 <= _zz_regVec_0_1;
          end
          if(_zz_2[1939]) begin
            regVec_1939 <= _zz_regVec_0_1;
          end
          if(_zz_2[1940]) begin
            regVec_1940 <= _zz_regVec_0_1;
          end
          if(_zz_2[1941]) begin
            regVec_1941 <= _zz_regVec_0_1;
          end
          if(_zz_2[1942]) begin
            regVec_1942 <= _zz_regVec_0_1;
          end
          if(_zz_2[1943]) begin
            regVec_1943 <= _zz_regVec_0_1;
          end
          if(_zz_2[1944]) begin
            regVec_1944 <= _zz_regVec_0_1;
          end
          if(_zz_2[1945]) begin
            regVec_1945 <= _zz_regVec_0_1;
          end
          if(_zz_2[1946]) begin
            regVec_1946 <= _zz_regVec_0_1;
          end
          if(_zz_2[1947]) begin
            regVec_1947 <= _zz_regVec_0_1;
          end
          if(_zz_2[1948]) begin
            regVec_1948 <= _zz_regVec_0_1;
          end
          if(_zz_2[1949]) begin
            regVec_1949 <= _zz_regVec_0_1;
          end
          if(_zz_2[1950]) begin
            regVec_1950 <= _zz_regVec_0_1;
          end
          if(_zz_2[1951]) begin
            regVec_1951 <= _zz_regVec_0_1;
          end
          if(_zz_2[1952]) begin
            regVec_1952 <= _zz_regVec_0_1;
          end
          if(_zz_2[1953]) begin
            regVec_1953 <= _zz_regVec_0_1;
          end
          if(_zz_2[1954]) begin
            regVec_1954 <= _zz_regVec_0_1;
          end
          if(_zz_2[1955]) begin
            regVec_1955 <= _zz_regVec_0_1;
          end
          if(_zz_2[1956]) begin
            regVec_1956 <= _zz_regVec_0_1;
          end
          if(_zz_2[1957]) begin
            regVec_1957 <= _zz_regVec_0_1;
          end
          if(_zz_2[1958]) begin
            regVec_1958 <= _zz_regVec_0_1;
          end
          if(_zz_2[1959]) begin
            regVec_1959 <= _zz_regVec_0_1;
          end
          if(_zz_2[1960]) begin
            regVec_1960 <= _zz_regVec_0_1;
          end
          if(_zz_2[1961]) begin
            regVec_1961 <= _zz_regVec_0_1;
          end
          if(_zz_2[1962]) begin
            regVec_1962 <= _zz_regVec_0_1;
          end
          if(_zz_2[1963]) begin
            regVec_1963 <= _zz_regVec_0_1;
          end
          if(_zz_2[1964]) begin
            regVec_1964 <= _zz_regVec_0_1;
          end
          if(_zz_2[1965]) begin
            regVec_1965 <= _zz_regVec_0_1;
          end
          if(_zz_2[1966]) begin
            regVec_1966 <= _zz_regVec_0_1;
          end
          if(_zz_2[1967]) begin
            regVec_1967 <= _zz_regVec_0_1;
          end
          if(_zz_2[1968]) begin
            regVec_1968 <= _zz_regVec_0_1;
          end
          if(_zz_2[1969]) begin
            regVec_1969 <= _zz_regVec_0_1;
          end
          if(_zz_2[1970]) begin
            regVec_1970 <= _zz_regVec_0_1;
          end
          if(_zz_2[1971]) begin
            regVec_1971 <= _zz_regVec_0_1;
          end
          if(_zz_2[1972]) begin
            regVec_1972 <= _zz_regVec_0_1;
          end
          if(_zz_2[1973]) begin
            regVec_1973 <= _zz_regVec_0_1;
          end
          if(_zz_2[1974]) begin
            regVec_1974 <= _zz_regVec_0_1;
          end
          if(_zz_2[1975]) begin
            regVec_1975 <= _zz_regVec_0_1;
          end
          if(_zz_2[1976]) begin
            regVec_1976 <= _zz_regVec_0_1;
          end
          if(_zz_2[1977]) begin
            regVec_1977 <= _zz_regVec_0_1;
          end
          if(_zz_2[1978]) begin
            regVec_1978 <= _zz_regVec_0_1;
          end
          if(_zz_2[1979]) begin
            regVec_1979 <= _zz_regVec_0_1;
          end
          if(_zz_2[1980]) begin
            regVec_1980 <= _zz_regVec_0_1;
          end
          if(_zz_2[1981]) begin
            regVec_1981 <= _zz_regVec_0_1;
          end
          if(_zz_2[1982]) begin
            regVec_1982 <= _zz_regVec_0_1;
          end
          if(_zz_2[1983]) begin
            regVec_1983 <= _zz_regVec_0_1;
          end
          if(_zz_2[1984]) begin
            regVec_1984 <= _zz_regVec_0_1;
          end
          if(_zz_2[1985]) begin
            regVec_1985 <= _zz_regVec_0_1;
          end
          if(_zz_2[1986]) begin
            regVec_1986 <= _zz_regVec_0_1;
          end
          if(_zz_2[1987]) begin
            regVec_1987 <= _zz_regVec_0_1;
          end
          if(_zz_2[1988]) begin
            regVec_1988 <= _zz_regVec_0_1;
          end
          if(_zz_2[1989]) begin
            regVec_1989 <= _zz_regVec_0_1;
          end
          if(_zz_2[1990]) begin
            regVec_1990 <= _zz_regVec_0_1;
          end
          if(_zz_2[1991]) begin
            regVec_1991 <= _zz_regVec_0_1;
          end
          if(_zz_2[1992]) begin
            regVec_1992 <= _zz_regVec_0_1;
          end
          if(_zz_2[1993]) begin
            regVec_1993 <= _zz_regVec_0_1;
          end
          if(_zz_2[1994]) begin
            regVec_1994 <= _zz_regVec_0_1;
          end
          if(_zz_2[1995]) begin
            regVec_1995 <= _zz_regVec_0_1;
          end
          if(_zz_2[1996]) begin
            regVec_1996 <= _zz_regVec_0_1;
          end
          if(_zz_2[1997]) begin
            regVec_1997 <= _zz_regVec_0_1;
          end
          if(_zz_2[1998]) begin
            regVec_1998 <= _zz_regVec_0_1;
          end
          if(_zz_2[1999]) begin
            regVec_1999 <= _zz_regVec_0_1;
          end
          if(_zz_2[2000]) begin
            regVec_2000 <= _zz_regVec_0_1;
          end
          if(_zz_2[2001]) begin
            regVec_2001 <= _zz_regVec_0_1;
          end
          if(_zz_2[2002]) begin
            regVec_2002 <= _zz_regVec_0_1;
          end
          if(_zz_2[2003]) begin
            regVec_2003 <= _zz_regVec_0_1;
          end
          if(_zz_2[2004]) begin
            regVec_2004 <= _zz_regVec_0_1;
          end
          if(_zz_2[2005]) begin
            regVec_2005 <= _zz_regVec_0_1;
          end
          if(_zz_2[2006]) begin
            regVec_2006 <= _zz_regVec_0_1;
          end
          if(_zz_2[2007]) begin
            regVec_2007 <= _zz_regVec_0_1;
          end
          if(_zz_2[2008]) begin
            regVec_2008 <= _zz_regVec_0_1;
          end
          if(_zz_2[2009]) begin
            regVec_2009 <= _zz_regVec_0_1;
          end
          if(_zz_2[2010]) begin
            regVec_2010 <= _zz_regVec_0_1;
          end
          if(_zz_2[2011]) begin
            regVec_2011 <= _zz_regVec_0_1;
          end
          if(_zz_2[2012]) begin
            regVec_2012 <= _zz_regVec_0_1;
          end
          if(_zz_2[2013]) begin
            regVec_2013 <= _zz_regVec_0_1;
          end
          if(_zz_2[2014]) begin
            regVec_2014 <= _zz_regVec_0_1;
          end
          if(_zz_2[2015]) begin
            regVec_2015 <= _zz_regVec_0_1;
          end
          if(_zz_2[2016]) begin
            regVec_2016 <= _zz_regVec_0_1;
          end
          if(_zz_2[2017]) begin
            regVec_2017 <= _zz_regVec_0_1;
          end
          if(_zz_2[2018]) begin
            regVec_2018 <= _zz_regVec_0_1;
          end
          if(_zz_2[2019]) begin
            regVec_2019 <= _zz_regVec_0_1;
          end
          if(_zz_2[2020]) begin
            regVec_2020 <= _zz_regVec_0_1;
          end
          if(_zz_2[2021]) begin
            regVec_2021 <= _zz_regVec_0_1;
          end
          if(_zz_2[2022]) begin
            regVec_2022 <= _zz_regVec_0_1;
          end
          if(_zz_2[2023]) begin
            regVec_2023 <= _zz_regVec_0_1;
          end
          if(_zz_2[2024]) begin
            regVec_2024 <= _zz_regVec_0_1;
          end
          if(_zz_2[2025]) begin
            regVec_2025 <= _zz_regVec_0_1;
          end
          if(_zz_2[2026]) begin
            regVec_2026 <= _zz_regVec_0_1;
          end
          if(_zz_2[2027]) begin
            regVec_2027 <= _zz_regVec_0_1;
          end
          if(_zz_2[2028]) begin
            regVec_2028 <= _zz_regVec_0_1;
          end
          if(_zz_2[2029]) begin
            regVec_2029 <= _zz_regVec_0_1;
          end
          if(_zz_2[2030]) begin
            regVec_2030 <= _zz_regVec_0_1;
          end
          if(_zz_2[2031]) begin
            regVec_2031 <= _zz_regVec_0_1;
          end
          if(_zz_2[2032]) begin
            regVec_2032 <= _zz_regVec_0_1;
          end
          if(_zz_2[2033]) begin
            regVec_2033 <= _zz_regVec_0_1;
          end
          if(_zz_2[2034]) begin
            regVec_2034 <= _zz_regVec_0_1;
          end
          if(_zz_2[2035]) begin
            regVec_2035 <= _zz_regVec_0_1;
          end
          if(_zz_2[2036]) begin
            regVec_2036 <= _zz_regVec_0_1;
          end
          if(_zz_2[2037]) begin
            regVec_2037 <= _zz_regVec_0_1;
          end
          if(_zz_2[2038]) begin
            regVec_2038 <= _zz_regVec_0_1;
          end
          if(_zz_2[2039]) begin
            regVec_2039 <= _zz_regVec_0_1;
          end
          if(_zz_2[2040]) begin
            regVec_2040 <= _zz_regVec_0_1;
          end
          if(_zz_2[2041]) begin
            regVec_2041 <= _zz_regVec_0_1;
          end
          if(_zz_2[2042]) begin
            regVec_2042 <= _zz_regVec_0_1;
          end
          if(_zz_2[2043]) begin
            regVec_2043 <= _zz_regVec_0_1;
          end
          if(_zz_2[2044]) begin
            regVec_2044 <= _zz_regVec_0_1;
          end
          if(_zz_2[2045]) begin
            regVec_2045 <= _zz_regVec_0_1;
          end
          if(_zz_2[2046]) begin
            regVec_2046 <= _zz_regVec_0_1;
          end
          if(_zz_2[2047]) begin
            regVec_2047 <= _zz_regVec_0_1;
          end
          if(_zz_2[2048]) begin
            regVec_2048 <= _zz_regVec_0_1;
          end
          if(_zz_2[2049]) begin
            regVec_2049 <= _zz_regVec_0_1;
          end
          if(_zz_2[2050]) begin
            regVec_2050 <= _zz_regVec_0_1;
          end
          if(_zz_2[2051]) begin
            regVec_2051 <= _zz_regVec_0_1;
          end
          if(_zz_2[2052]) begin
            regVec_2052 <= _zz_regVec_0_1;
          end
          if(_zz_2[2053]) begin
            regVec_2053 <= _zz_regVec_0_1;
          end
          if(_zz_2[2054]) begin
            regVec_2054 <= _zz_regVec_0_1;
          end
          if(_zz_2[2055]) begin
            regVec_2055 <= _zz_regVec_0_1;
          end
          if(_zz_2[2056]) begin
            regVec_2056 <= _zz_regVec_0_1;
          end
          if(_zz_2[2057]) begin
            regVec_2057 <= _zz_regVec_0_1;
          end
          if(_zz_2[2058]) begin
            regVec_2058 <= _zz_regVec_0_1;
          end
          if(_zz_2[2059]) begin
            regVec_2059 <= _zz_regVec_0_1;
          end
          if(_zz_2[2060]) begin
            regVec_2060 <= _zz_regVec_0_1;
          end
          if(_zz_2[2061]) begin
            regVec_2061 <= _zz_regVec_0_1;
          end
          if(_zz_2[2062]) begin
            regVec_2062 <= _zz_regVec_0_1;
          end
          if(_zz_2[2063]) begin
            regVec_2063 <= _zz_regVec_0_1;
          end
          if(_zz_2[2064]) begin
            regVec_2064 <= _zz_regVec_0_1;
          end
          if(_zz_2[2065]) begin
            regVec_2065 <= _zz_regVec_0_1;
          end
          if(_zz_2[2066]) begin
            regVec_2066 <= _zz_regVec_0_1;
          end
          if(_zz_2[2067]) begin
            regVec_2067 <= _zz_regVec_0_1;
          end
          if(_zz_2[2068]) begin
            regVec_2068 <= _zz_regVec_0_1;
          end
          if(_zz_2[2069]) begin
            regVec_2069 <= _zz_regVec_0_1;
          end
          if(_zz_2[2070]) begin
            regVec_2070 <= _zz_regVec_0_1;
          end
          if(_zz_2[2071]) begin
            regVec_2071 <= _zz_regVec_0_1;
          end
          if(_zz_2[2072]) begin
            regVec_2072 <= _zz_regVec_0_1;
          end
          if(_zz_2[2073]) begin
            regVec_2073 <= _zz_regVec_0_1;
          end
          if(_zz_2[2074]) begin
            regVec_2074 <= _zz_regVec_0_1;
          end
          if(_zz_2[2075]) begin
            regVec_2075 <= _zz_regVec_0_1;
          end
          if(_zz_2[2076]) begin
            regVec_2076 <= _zz_regVec_0_1;
          end
          if(_zz_2[2077]) begin
            regVec_2077 <= _zz_regVec_0_1;
          end
          if(_zz_2[2078]) begin
            regVec_2078 <= _zz_regVec_0_1;
          end
          if(_zz_2[2079]) begin
            regVec_2079 <= _zz_regVec_0_1;
          end
          if(_zz_2[2080]) begin
            regVec_2080 <= _zz_regVec_0_1;
          end
          if(_zz_2[2081]) begin
            regVec_2081 <= _zz_regVec_0_1;
          end
          if(_zz_2[2082]) begin
            regVec_2082 <= _zz_regVec_0_1;
          end
          if(_zz_2[2083]) begin
            regVec_2083 <= _zz_regVec_0_1;
          end
          if(_zz_2[2084]) begin
            regVec_2084 <= _zz_regVec_0_1;
          end
          if(_zz_2[2085]) begin
            regVec_2085 <= _zz_regVec_0_1;
          end
          if(_zz_2[2086]) begin
            regVec_2086 <= _zz_regVec_0_1;
          end
          if(_zz_2[2087]) begin
            regVec_2087 <= _zz_regVec_0_1;
          end
          if(_zz_2[2088]) begin
            regVec_2088 <= _zz_regVec_0_1;
          end
          if(_zz_2[2089]) begin
            regVec_2089 <= _zz_regVec_0_1;
          end
          if(_zz_2[2090]) begin
            regVec_2090 <= _zz_regVec_0_1;
          end
          if(_zz_2[2091]) begin
            regVec_2091 <= _zz_regVec_0_1;
          end
          if(_zz_2[2092]) begin
            regVec_2092 <= _zz_regVec_0_1;
          end
          if(_zz_2[2093]) begin
            regVec_2093 <= _zz_regVec_0_1;
          end
          if(_zz_2[2094]) begin
            regVec_2094 <= _zz_regVec_0_1;
          end
          if(_zz_2[2095]) begin
            regVec_2095 <= _zz_regVec_0_1;
          end
          if(_zz_2[2096]) begin
            regVec_2096 <= _zz_regVec_0_1;
          end
          if(_zz_2[2097]) begin
            regVec_2097 <= _zz_regVec_0_1;
          end
          if(_zz_2[2098]) begin
            regVec_2098 <= _zz_regVec_0_1;
          end
          if(_zz_2[2099]) begin
            regVec_2099 <= _zz_regVec_0_1;
          end
          if(_zz_2[2100]) begin
            regVec_2100 <= _zz_regVec_0_1;
          end
          if(_zz_2[2101]) begin
            regVec_2101 <= _zz_regVec_0_1;
          end
          if(_zz_2[2102]) begin
            regVec_2102 <= _zz_regVec_0_1;
          end
          if(_zz_2[2103]) begin
            regVec_2103 <= _zz_regVec_0_1;
          end
          if(_zz_2[2104]) begin
            regVec_2104 <= _zz_regVec_0_1;
          end
          if(_zz_2[2105]) begin
            regVec_2105 <= _zz_regVec_0_1;
          end
          if(_zz_2[2106]) begin
            regVec_2106 <= _zz_regVec_0_1;
          end
          if(_zz_2[2107]) begin
            regVec_2107 <= _zz_regVec_0_1;
          end
          if(_zz_2[2108]) begin
            regVec_2108 <= _zz_regVec_0_1;
          end
          if(_zz_2[2109]) begin
            regVec_2109 <= _zz_regVec_0_1;
          end
          if(_zz_2[2110]) begin
            regVec_2110 <= _zz_regVec_0_1;
          end
          if(_zz_2[2111]) begin
            regVec_2111 <= _zz_regVec_0_1;
          end
          if(_zz_2[2112]) begin
            regVec_2112 <= _zz_regVec_0_1;
          end
          if(_zz_2[2113]) begin
            regVec_2113 <= _zz_regVec_0_1;
          end
          if(_zz_2[2114]) begin
            regVec_2114 <= _zz_regVec_0_1;
          end
          if(_zz_2[2115]) begin
            regVec_2115 <= _zz_regVec_0_1;
          end
          if(_zz_2[2116]) begin
            regVec_2116 <= _zz_regVec_0_1;
          end
          if(_zz_2[2117]) begin
            regVec_2117 <= _zz_regVec_0_1;
          end
          if(_zz_2[2118]) begin
            regVec_2118 <= _zz_regVec_0_1;
          end
          if(_zz_2[2119]) begin
            regVec_2119 <= _zz_regVec_0_1;
          end
          if(_zz_2[2120]) begin
            regVec_2120 <= _zz_regVec_0_1;
          end
          if(_zz_2[2121]) begin
            regVec_2121 <= _zz_regVec_0_1;
          end
          if(_zz_2[2122]) begin
            regVec_2122 <= _zz_regVec_0_1;
          end
          if(_zz_2[2123]) begin
            regVec_2123 <= _zz_regVec_0_1;
          end
          if(_zz_2[2124]) begin
            regVec_2124 <= _zz_regVec_0_1;
          end
          if(_zz_2[2125]) begin
            regVec_2125 <= _zz_regVec_0_1;
          end
          if(_zz_2[2126]) begin
            regVec_2126 <= _zz_regVec_0_1;
          end
          if(_zz_2[2127]) begin
            regVec_2127 <= _zz_regVec_0_1;
          end
          if(_zz_2[2128]) begin
            regVec_2128 <= _zz_regVec_0_1;
          end
          if(_zz_2[2129]) begin
            regVec_2129 <= _zz_regVec_0_1;
          end
          if(_zz_2[2130]) begin
            regVec_2130 <= _zz_regVec_0_1;
          end
          if(_zz_2[2131]) begin
            regVec_2131 <= _zz_regVec_0_1;
          end
          if(_zz_2[2132]) begin
            regVec_2132 <= _zz_regVec_0_1;
          end
          if(_zz_2[2133]) begin
            regVec_2133 <= _zz_regVec_0_1;
          end
          if(_zz_2[2134]) begin
            regVec_2134 <= _zz_regVec_0_1;
          end
          if(_zz_2[2135]) begin
            regVec_2135 <= _zz_regVec_0_1;
          end
          if(_zz_2[2136]) begin
            regVec_2136 <= _zz_regVec_0_1;
          end
          if(_zz_2[2137]) begin
            regVec_2137 <= _zz_regVec_0_1;
          end
          if(_zz_2[2138]) begin
            regVec_2138 <= _zz_regVec_0_1;
          end
          if(_zz_2[2139]) begin
            regVec_2139 <= _zz_regVec_0_1;
          end
          if(_zz_2[2140]) begin
            regVec_2140 <= _zz_regVec_0_1;
          end
          if(_zz_2[2141]) begin
            regVec_2141 <= _zz_regVec_0_1;
          end
          if(_zz_2[2142]) begin
            regVec_2142 <= _zz_regVec_0_1;
          end
          if(_zz_2[2143]) begin
            regVec_2143 <= _zz_regVec_0_1;
          end
          if(_zz_2[2144]) begin
            regVec_2144 <= _zz_regVec_0_1;
          end
          if(_zz_2[2145]) begin
            regVec_2145 <= _zz_regVec_0_1;
          end
          if(_zz_2[2146]) begin
            regVec_2146 <= _zz_regVec_0_1;
          end
          if(_zz_2[2147]) begin
            regVec_2147 <= _zz_regVec_0_1;
          end
          if(_zz_2[2148]) begin
            regVec_2148 <= _zz_regVec_0_1;
          end
          if(_zz_2[2149]) begin
            regVec_2149 <= _zz_regVec_0_1;
          end
          if(_zz_2[2150]) begin
            regVec_2150 <= _zz_regVec_0_1;
          end
          if(_zz_2[2151]) begin
            regVec_2151 <= _zz_regVec_0_1;
          end
          if(_zz_2[2152]) begin
            regVec_2152 <= _zz_regVec_0_1;
          end
          if(_zz_2[2153]) begin
            regVec_2153 <= _zz_regVec_0_1;
          end
          if(_zz_2[2154]) begin
            regVec_2154 <= _zz_regVec_0_1;
          end
          if(_zz_2[2155]) begin
            regVec_2155 <= _zz_regVec_0_1;
          end
          if(_zz_2[2156]) begin
            regVec_2156 <= _zz_regVec_0_1;
          end
          if(_zz_2[2157]) begin
            regVec_2157 <= _zz_regVec_0_1;
          end
          if(_zz_2[2158]) begin
            regVec_2158 <= _zz_regVec_0_1;
          end
          if(_zz_2[2159]) begin
            regVec_2159 <= _zz_regVec_0_1;
          end
          if(_zz_2[2160]) begin
            regVec_2160 <= _zz_regVec_0_1;
          end
          if(_zz_2[2161]) begin
            regVec_2161 <= _zz_regVec_0_1;
          end
          if(_zz_2[2162]) begin
            regVec_2162 <= _zz_regVec_0_1;
          end
          if(_zz_2[2163]) begin
            regVec_2163 <= _zz_regVec_0_1;
          end
          if(_zz_2[2164]) begin
            regVec_2164 <= _zz_regVec_0_1;
          end
          if(_zz_2[2165]) begin
            regVec_2165 <= _zz_regVec_0_1;
          end
          if(_zz_2[2166]) begin
            regVec_2166 <= _zz_regVec_0_1;
          end
          if(_zz_2[2167]) begin
            regVec_2167 <= _zz_regVec_0_1;
          end
          if(_zz_2[2168]) begin
            regVec_2168 <= _zz_regVec_0_1;
          end
          if(_zz_2[2169]) begin
            regVec_2169 <= _zz_regVec_0_1;
          end
          if(_zz_2[2170]) begin
            regVec_2170 <= _zz_regVec_0_1;
          end
          if(_zz_2[2171]) begin
            regVec_2171 <= _zz_regVec_0_1;
          end
          if(_zz_2[2172]) begin
            regVec_2172 <= _zz_regVec_0_1;
          end
          if(_zz_2[2173]) begin
            regVec_2173 <= _zz_regVec_0_1;
          end
          if(_zz_2[2174]) begin
            regVec_2174 <= _zz_regVec_0_1;
          end
          if(_zz_2[2175]) begin
            regVec_2175 <= _zz_regVec_0_1;
          end
          if(_zz_2[2176]) begin
            regVec_2176 <= _zz_regVec_0_1;
          end
          if(_zz_2[2177]) begin
            regVec_2177 <= _zz_regVec_0_1;
          end
          if(_zz_2[2178]) begin
            regVec_2178 <= _zz_regVec_0_1;
          end
          if(_zz_2[2179]) begin
            regVec_2179 <= _zz_regVec_0_1;
          end
          if(_zz_2[2180]) begin
            regVec_2180 <= _zz_regVec_0_1;
          end
          if(_zz_2[2181]) begin
            regVec_2181 <= _zz_regVec_0_1;
          end
          if(_zz_2[2182]) begin
            regVec_2182 <= _zz_regVec_0_1;
          end
          if(_zz_2[2183]) begin
            regVec_2183 <= _zz_regVec_0_1;
          end
          if(_zz_2[2184]) begin
            regVec_2184 <= _zz_regVec_0_1;
          end
          if(_zz_2[2185]) begin
            regVec_2185 <= _zz_regVec_0_1;
          end
          if(_zz_2[2186]) begin
            regVec_2186 <= _zz_regVec_0_1;
          end
          if(_zz_2[2187]) begin
            regVec_2187 <= _zz_regVec_0_1;
          end
          if(_zz_2[2188]) begin
            regVec_2188 <= _zz_regVec_0_1;
          end
          if(_zz_2[2189]) begin
            regVec_2189 <= _zz_regVec_0_1;
          end
          if(_zz_2[2190]) begin
            regVec_2190 <= _zz_regVec_0_1;
          end
          if(_zz_2[2191]) begin
            regVec_2191 <= _zz_regVec_0_1;
          end
          if(_zz_2[2192]) begin
            regVec_2192 <= _zz_regVec_0_1;
          end
          if(_zz_2[2193]) begin
            regVec_2193 <= _zz_regVec_0_1;
          end
          if(_zz_2[2194]) begin
            regVec_2194 <= _zz_regVec_0_1;
          end
          if(_zz_2[2195]) begin
            regVec_2195 <= _zz_regVec_0_1;
          end
          if(_zz_2[2196]) begin
            regVec_2196 <= _zz_regVec_0_1;
          end
          if(_zz_2[2197]) begin
            regVec_2197 <= _zz_regVec_0_1;
          end
          if(_zz_2[2198]) begin
            regVec_2198 <= _zz_regVec_0_1;
          end
          if(_zz_2[2199]) begin
            regVec_2199 <= _zz_regVec_0_1;
          end
          if(_zz_2[2200]) begin
            regVec_2200 <= _zz_regVec_0_1;
          end
          if(_zz_2[2201]) begin
            regVec_2201 <= _zz_regVec_0_1;
          end
          if(_zz_2[2202]) begin
            regVec_2202 <= _zz_regVec_0_1;
          end
          if(_zz_2[2203]) begin
            regVec_2203 <= _zz_regVec_0_1;
          end
          if(_zz_2[2204]) begin
            regVec_2204 <= _zz_regVec_0_1;
          end
          if(_zz_2[2205]) begin
            regVec_2205 <= _zz_regVec_0_1;
          end
          if(_zz_2[2206]) begin
            regVec_2206 <= _zz_regVec_0_1;
          end
          if(_zz_2[2207]) begin
            regVec_2207 <= _zz_regVec_0_1;
          end
          if(_zz_2[2208]) begin
            regVec_2208 <= _zz_regVec_0_1;
          end
          if(_zz_2[2209]) begin
            regVec_2209 <= _zz_regVec_0_1;
          end
          if(_zz_2[2210]) begin
            regVec_2210 <= _zz_regVec_0_1;
          end
          if(_zz_2[2211]) begin
            regVec_2211 <= _zz_regVec_0_1;
          end
          if(_zz_2[2212]) begin
            regVec_2212 <= _zz_regVec_0_1;
          end
          if(_zz_2[2213]) begin
            regVec_2213 <= _zz_regVec_0_1;
          end
          if(_zz_2[2214]) begin
            regVec_2214 <= _zz_regVec_0_1;
          end
          if(_zz_2[2215]) begin
            regVec_2215 <= _zz_regVec_0_1;
          end
          if(_zz_2[2216]) begin
            regVec_2216 <= _zz_regVec_0_1;
          end
          if(_zz_2[2217]) begin
            regVec_2217 <= _zz_regVec_0_1;
          end
          if(_zz_2[2218]) begin
            regVec_2218 <= _zz_regVec_0_1;
          end
          if(_zz_2[2219]) begin
            regVec_2219 <= _zz_regVec_0_1;
          end
          if(_zz_2[2220]) begin
            regVec_2220 <= _zz_regVec_0_1;
          end
          if(_zz_2[2221]) begin
            regVec_2221 <= _zz_regVec_0_1;
          end
          if(_zz_2[2222]) begin
            regVec_2222 <= _zz_regVec_0_1;
          end
          if(_zz_2[2223]) begin
            regVec_2223 <= _zz_regVec_0_1;
          end
          if(_zz_2[2224]) begin
            regVec_2224 <= _zz_regVec_0_1;
          end
          if(_zz_2[2225]) begin
            regVec_2225 <= _zz_regVec_0_1;
          end
          if(_zz_2[2226]) begin
            regVec_2226 <= _zz_regVec_0_1;
          end
          if(_zz_2[2227]) begin
            regVec_2227 <= _zz_regVec_0_1;
          end
          if(_zz_2[2228]) begin
            regVec_2228 <= _zz_regVec_0_1;
          end
          if(_zz_2[2229]) begin
            regVec_2229 <= _zz_regVec_0_1;
          end
          if(_zz_2[2230]) begin
            regVec_2230 <= _zz_regVec_0_1;
          end
          if(_zz_2[2231]) begin
            regVec_2231 <= _zz_regVec_0_1;
          end
          if(_zz_2[2232]) begin
            regVec_2232 <= _zz_regVec_0_1;
          end
          if(_zz_2[2233]) begin
            regVec_2233 <= _zz_regVec_0_1;
          end
          if(_zz_2[2234]) begin
            regVec_2234 <= _zz_regVec_0_1;
          end
          if(_zz_2[2235]) begin
            regVec_2235 <= _zz_regVec_0_1;
          end
          if(_zz_2[2236]) begin
            regVec_2236 <= _zz_regVec_0_1;
          end
          if(_zz_2[2237]) begin
            regVec_2237 <= _zz_regVec_0_1;
          end
          if(_zz_2[2238]) begin
            regVec_2238 <= _zz_regVec_0_1;
          end
          if(_zz_2[2239]) begin
            regVec_2239 <= _zz_regVec_0_1;
          end
          if(_zz_2[2240]) begin
            regVec_2240 <= _zz_regVec_0_1;
          end
          if(_zz_2[2241]) begin
            regVec_2241 <= _zz_regVec_0_1;
          end
          if(_zz_2[2242]) begin
            regVec_2242 <= _zz_regVec_0_1;
          end
          if(_zz_2[2243]) begin
            regVec_2243 <= _zz_regVec_0_1;
          end
          if(_zz_2[2244]) begin
            regVec_2244 <= _zz_regVec_0_1;
          end
          if(_zz_2[2245]) begin
            regVec_2245 <= _zz_regVec_0_1;
          end
          if(_zz_2[2246]) begin
            regVec_2246 <= _zz_regVec_0_1;
          end
          if(_zz_2[2247]) begin
            regVec_2247 <= _zz_regVec_0_1;
          end
          if(_zz_2[2248]) begin
            regVec_2248 <= _zz_regVec_0_1;
          end
          if(_zz_2[2249]) begin
            regVec_2249 <= _zz_regVec_0_1;
          end
          if(_zz_2[2250]) begin
            regVec_2250 <= _zz_regVec_0_1;
          end
          if(_zz_2[2251]) begin
            regVec_2251 <= _zz_regVec_0_1;
          end
          if(_zz_2[2252]) begin
            regVec_2252 <= _zz_regVec_0_1;
          end
          if(_zz_2[2253]) begin
            regVec_2253 <= _zz_regVec_0_1;
          end
          if(_zz_2[2254]) begin
            regVec_2254 <= _zz_regVec_0_1;
          end
          if(_zz_2[2255]) begin
            regVec_2255 <= _zz_regVec_0_1;
          end
          if(_zz_2[2256]) begin
            regVec_2256 <= _zz_regVec_0_1;
          end
          if(_zz_2[2257]) begin
            regVec_2257 <= _zz_regVec_0_1;
          end
          if(_zz_2[2258]) begin
            regVec_2258 <= _zz_regVec_0_1;
          end
          if(_zz_2[2259]) begin
            regVec_2259 <= _zz_regVec_0_1;
          end
          if(_zz_2[2260]) begin
            regVec_2260 <= _zz_regVec_0_1;
          end
          if(_zz_2[2261]) begin
            regVec_2261 <= _zz_regVec_0_1;
          end
          if(_zz_2[2262]) begin
            regVec_2262 <= _zz_regVec_0_1;
          end
          if(_zz_2[2263]) begin
            regVec_2263 <= _zz_regVec_0_1;
          end
          if(_zz_2[2264]) begin
            regVec_2264 <= _zz_regVec_0_1;
          end
          if(_zz_2[2265]) begin
            regVec_2265 <= _zz_regVec_0_1;
          end
          if(_zz_2[2266]) begin
            regVec_2266 <= _zz_regVec_0_1;
          end
          if(_zz_2[2267]) begin
            regVec_2267 <= _zz_regVec_0_1;
          end
          if(_zz_2[2268]) begin
            regVec_2268 <= _zz_regVec_0_1;
          end
          if(_zz_2[2269]) begin
            regVec_2269 <= _zz_regVec_0_1;
          end
          if(_zz_2[2270]) begin
            regVec_2270 <= _zz_regVec_0_1;
          end
          if(_zz_2[2271]) begin
            regVec_2271 <= _zz_regVec_0_1;
          end
          if(_zz_2[2272]) begin
            regVec_2272 <= _zz_regVec_0_1;
          end
          if(_zz_2[2273]) begin
            regVec_2273 <= _zz_regVec_0_1;
          end
          if(_zz_2[2274]) begin
            regVec_2274 <= _zz_regVec_0_1;
          end
          if(_zz_2[2275]) begin
            regVec_2275 <= _zz_regVec_0_1;
          end
          if(_zz_2[2276]) begin
            regVec_2276 <= _zz_regVec_0_1;
          end
          if(_zz_2[2277]) begin
            regVec_2277 <= _zz_regVec_0_1;
          end
          if(_zz_2[2278]) begin
            regVec_2278 <= _zz_regVec_0_1;
          end
          if(_zz_2[2279]) begin
            regVec_2279 <= _zz_regVec_0_1;
          end
          if(_zz_2[2280]) begin
            regVec_2280 <= _zz_regVec_0_1;
          end
          if(_zz_2[2281]) begin
            regVec_2281 <= _zz_regVec_0_1;
          end
          if(_zz_2[2282]) begin
            regVec_2282 <= _zz_regVec_0_1;
          end
          if(_zz_2[2283]) begin
            regVec_2283 <= _zz_regVec_0_1;
          end
          if(_zz_2[2284]) begin
            regVec_2284 <= _zz_regVec_0_1;
          end
          if(_zz_2[2285]) begin
            regVec_2285 <= _zz_regVec_0_1;
          end
          if(_zz_2[2286]) begin
            regVec_2286 <= _zz_regVec_0_1;
          end
          if(_zz_2[2287]) begin
            regVec_2287 <= _zz_regVec_0_1;
          end
          if(_zz_2[2288]) begin
            regVec_2288 <= _zz_regVec_0_1;
          end
          if(_zz_2[2289]) begin
            regVec_2289 <= _zz_regVec_0_1;
          end
          if(_zz_2[2290]) begin
            regVec_2290 <= _zz_regVec_0_1;
          end
          if(_zz_2[2291]) begin
            regVec_2291 <= _zz_regVec_0_1;
          end
          if(_zz_2[2292]) begin
            regVec_2292 <= _zz_regVec_0_1;
          end
          if(_zz_2[2293]) begin
            regVec_2293 <= _zz_regVec_0_1;
          end
          if(_zz_2[2294]) begin
            regVec_2294 <= _zz_regVec_0_1;
          end
          if(_zz_2[2295]) begin
            regVec_2295 <= _zz_regVec_0_1;
          end
          if(_zz_2[2296]) begin
            regVec_2296 <= _zz_regVec_0_1;
          end
          if(_zz_2[2297]) begin
            regVec_2297 <= _zz_regVec_0_1;
          end
          if(_zz_2[2298]) begin
            regVec_2298 <= _zz_regVec_0_1;
          end
          if(_zz_2[2299]) begin
            regVec_2299 <= _zz_regVec_0_1;
          end
          if(_zz_2[2300]) begin
            regVec_2300 <= _zz_regVec_0_1;
          end
          if(_zz_2[2301]) begin
            regVec_2301 <= _zz_regVec_0_1;
          end
          if(_zz_2[2302]) begin
            regVec_2302 <= _zz_regVec_0_1;
          end
          if(_zz_2[2303]) begin
            regVec_2303 <= _zz_regVec_0_1;
          end
          if(_zz_2[2304]) begin
            regVec_2304 <= _zz_regVec_0_1;
          end
          if(_zz_2[2305]) begin
            regVec_2305 <= _zz_regVec_0_1;
          end
          if(_zz_2[2306]) begin
            regVec_2306 <= _zz_regVec_0_1;
          end
          if(_zz_2[2307]) begin
            regVec_2307 <= _zz_regVec_0_1;
          end
          if(_zz_2[2308]) begin
            regVec_2308 <= _zz_regVec_0_1;
          end
          if(_zz_2[2309]) begin
            regVec_2309 <= _zz_regVec_0_1;
          end
          if(_zz_2[2310]) begin
            regVec_2310 <= _zz_regVec_0_1;
          end
          if(_zz_2[2311]) begin
            regVec_2311 <= _zz_regVec_0_1;
          end
          if(_zz_2[2312]) begin
            regVec_2312 <= _zz_regVec_0_1;
          end
          if(_zz_2[2313]) begin
            regVec_2313 <= _zz_regVec_0_1;
          end
          if(_zz_2[2314]) begin
            regVec_2314 <= _zz_regVec_0_1;
          end
          if(_zz_2[2315]) begin
            regVec_2315 <= _zz_regVec_0_1;
          end
          if(_zz_2[2316]) begin
            regVec_2316 <= _zz_regVec_0_1;
          end
          if(_zz_2[2317]) begin
            regVec_2317 <= _zz_regVec_0_1;
          end
          if(_zz_2[2318]) begin
            regVec_2318 <= _zz_regVec_0_1;
          end
          if(_zz_2[2319]) begin
            regVec_2319 <= _zz_regVec_0_1;
          end
          if(_zz_2[2320]) begin
            regVec_2320 <= _zz_regVec_0_1;
          end
          if(_zz_2[2321]) begin
            regVec_2321 <= _zz_regVec_0_1;
          end
          if(_zz_2[2322]) begin
            regVec_2322 <= _zz_regVec_0_1;
          end
          if(_zz_2[2323]) begin
            regVec_2323 <= _zz_regVec_0_1;
          end
          if(_zz_2[2324]) begin
            regVec_2324 <= _zz_regVec_0_1;
          end
          if(_zz_2[2325]) begin
            regVec_2325 <= _zz_regVec_0_1;
          end
          if(_zz_2[2326]) begin
            regVec_2326 <= _zz_regVec_0_1;
          end
          if(_zz_2[2327]) begin
            regVec_2327 <= _zz_regVec_0_1;
          end
          if(_zz_2[2328]) begin
            regVec_2328 <= _zz_regVec_0_1;
          end
          if(_zz_2[2329]) begin
            regVec_2329 <= _zz_regVec_0_1;
          end
          if(_zz_2[2330]) begin
            regVec_2330 <= _zz_regVec_0_1;
          end
          if(_zz_2[2331]) begin
            regVec_2331 <= _zz_regVec_0_1;
          end
          if(_zz_2[2332]) begin
            regVec_2332 <= _zz_regVec_0_1;
          end
          if(_zz_2[2333]) begin
            regVec_2333 <= _zz_regVec_0_1;
          end
          if(_zz_2[2334]) begin
            regVec_2334 <= _zz_regVec_0_1;
          end
          if(_zz_2[2335]) begin
            regVec_2335 <= _zz_regVec_0_1;
          end
          if(_zz_2[2336]) begin
            regVec_2336 <= _zz_regVec_0_1;
          end
          if(_zz_2[2337]) begin
            regVec_2337 <= _zz_regVec_0_1;
          end
          if(_zz_2[2338]) begin
            regVec_2338 <= _zz_regVec_0_1;
          end
          if(_zz_2[2339]) begin
            regVec_2339 <= _zz_regVec_0_1;
          end
          if(_zz_2[2340]) begin
            regVec_2340 <= _zz_regVec_0_1;
          end
          if(_zz_2[2341]) begin
            regVec_2341 <= _zz_regVec_0_1;
          end
          if(_zz_2[2342]) begin
            regVec_2342 <= _zz_regVec_0_1;
          end
          if(_zz_2[2343]) begin
            regVec_2343 <= _zz_regVec_0_1;
          end
          if(_zz_2[2344]) begin
            regVec_2344 <= _zz_regVec_0_1;
          end
          if(_zz_2[2345]) begin
            regVec_2345 <= _zz_regVec_0_1;
          end
          if(_zz_2[2346]) begin
            regVec_2346 <= _zz_regVec_0_1;
          end
          if(_zz_2[2347]) begin
            regVec_2347 <= _zz_regVec_0_1;
          end
          if(_zz_2[2348]) begin
            regVec_2348 <= _zz_regVec_0_1;
          end
          if(_zz_2[2349]) begin
            regVec_2349 <= _zz_regVec_0_1;
          end
          if(_zz_2[2350]) begin
            regVec_2350 <= _zz_regVec_0_1;
          end
          if(_zz_2[2351]) begin
            regVec_2351 <= _zz_regVec_0_1;
          end
          if(_zz_2[2352]) begin
            regVec_2352 <= _zz_regVec_0_1;
          end
          if(_zz_2[2353]) begin
            regVec_2353 <= _zz_regVec_0_1;
          end
          if(_zz_2[2354]) begin
            regVec_2354 <= _zz_regVec_0_1;
          end
          if(_zz_2[2355]) begin
            regVec_2355 <= _zz_regVec_0_1;
          end
          if(_zz_2[2356]) begin
            regVec_2356 <= _zz_regVec_0_1;
          end
          if(_zz_2[2357]) begin
            regVec_2357 <= _zz_regVec_0_1;
          end
          if(_zz_2[2358]) begin
            regVec_2358 <= _zz_regVec_0_1;
          end
          if(_zz_2[2359]) begin
            regVec_2359 <= _zz_regVec_0_1;
          end
          if(_zz_2[2360]) begin
            regVec_2360 <= _zz_regVec_0_1;
          end
          if(_zz_2[2361]) begin
            regVec_2361 <= _zz_regVec_0_1;
          end
          if(_zz_2[2362]) begin
            regVec_2362 <= _zz_regVec_0_1;
          end
          if(_zz_2[2363]) begin
            regVec_2363 <= _zz_regVec_0_1;
          end
          if(_zz_2[2364]) begin
            regVec_2364 <= _zz_regVec_0_1;
          end
          if(_zz_2[2365]) begin
            regVec_2365 <= _zz_regVec_0_1;
          end
          if(_zz_2[2366]) begin
            regVec_2366 <= _zz_regVec_0_1;
          end
          if(_zz_2[2367]) begin
            regVec_2367 <= _zz_regVec_0_1;
          end
          if(_zz_2[2368]) begin
            regVec_2368 <= _zz_regVec_0_1;
          end
          if(_zz_2[2369]) begin
            regVec_2369 <= _zz_regVec_0_1;
          end
          if(_zz_2[2370]) begin
            regVec_2370 <= _zz_regVec_0_1;
          end
          if(_zz_2[2371]) begin
            regVec_2371 <= _zz_regVec_0_1;
          end
          if(_zz_2[2372]) begin
            regVec_2372 <= _zz_regVec_0_1;
          end
          if(_zz_2[2373]) begin
            regVec_2373 <= _zz_regVec_0_1;
          end
          if(_zz_2[2374]) begin
            regVec_2374 <= _zz_regVec_0_1;
          end
          if(_zz_2[2375]) begin
            regVec_2375 <= _zz_regVec_0_1;
          end
          if(_zz_2[2376]) begin
            regVec_2376 <= _zz_regVec_0_1;
          end
          if(_zz_2[2377]) begin
            regVec_2377 <= _zz_regVec_0_1;
          end
          if(_zz_2[2378]) begin
            regVec_2378 <= _zz_regVec_0_1;
          end
          if(_zz_2[2379]) begin
            regVec_2379 <= _zz_regVec_0_1;
          end
          if(_zz_2[2380]) begin
            regVec_2380 <= _zz_regVec_0_1;
          end
          if(_zz_2[2381]) begin
            regVec_2381 <= _zz_regVec_0_1;
          end
          if(_zz_2[2382]) begin
            regVec_2382 <= _zz_regVec_0_1;
          end
          if(_zz_2[2383]) begin
            regVec_2383 <= _zz_regVec_0_1;
          end
          if(_zz_2[2384]) begin
            regVec_2384 <= _zz_regVec_0_1;
          end
          if(_zz_2[2385]) begin
            regVec_2385 <= _zz_regVec_0_1;
          end
          if(_zz_2[2386]) begin
            regVec_2386 <= _zz_regVec_0_1;
          end
          if(_zz_2[2387]) begin
            regVec_2387 <= _zz_regVec_0_1;
          end
          if(_zz_2[2388]) begin
            regVec_2388 <= _zz_regVec_0_1;
          end
          if(_zz_2[2389]) begin
            regVec_2389 <= _zz_regVec_0_1;
          end
          if(_zz_2[2390]) begin
            regVec_2390 <= _zz_regVec_0_1;
          end
          if(_zz_2[2391]) begin
            regVec_2391 <= _zz_regVec_0_1;
          end
          if(_zz_2[2392]) begin
            regVec_2392 <= _zz_regVec_0_1;
          end
          if(_zz_2[2393]) begin
            regVec_2393 <= _zz_regVec_0_1;
          end
          if(_zz_2[2394]) begin
            regVec_2394 <= _zz_regVec_0_1;
          end
          if(_zz_2[2395]) begin
            regVec_2395 <= _zz_regVec_0_1;
          end
          if(_zz_2[2396]) begin
            regVec_2396 <= _zz_regVec_0_1;
          end
          if(_zz_2[2397]) begin
            regVec_2397 <= _zz_regVec_0_1;
          end
          if(_zz_2[2398]) begin
            regVec_2398 <= _zz_regVec_0_1;
          end
          if(_zz_2[2399]) begin
            regVec_2399 <= _zz_regVec_0_1;
          end
          if(_zz_2[2400]) begin
            regVec_2400 <= _zz_regVec_0_1;
          end
          if(_zz_2[2401]) begin
            regVec_2401 <= _zz_regVec_0_1;
          end
          if(_zz_2[2402]) begin
            regVec_2402 <= _zz_regVec_0_1;
          end
          if(_zz_2[2403]) begin
            regVec_2403 <= _zz_regVec_0_1;
          end
          if(_zz_2[2404]) begin
            regVec_2404 <= _zz_regVec_0_1;
          end
          if(_zz_2[2405]) begin
            regVec_2405 <= _zz_regVec_0_1;
          end
          if(_zz_2[2406]) begin
            regVec_2406 <= _zz_regVec_0_1;
          end
          if(_zz_2[2407]) begin
            regVec_2407 <= _zz_regVec_0_1;
          end
          if(_zz_2[2408]) begin
            regVec_2408 <= _zz_regVec_0_1;
          end
          if(_zz_2[2409]) begin
            regVec_2409 <= _zz_regVec_0_1;
          end
          if(_zz_2[2410]) begin
            regVec_2410 <= _zz_regVec_0_1;
          end
          if(_zz_2[2411]) begin
            regVec_2411 <= _zz_regVec_0_1;
          end
          if(_zz_2[2412]) begin
            regVec_2412 <= _zz_regVec_0_1;
          end
          if(_zz_2[2413]) begin
            regVec_2413 <= _zz_regVec_0_1;
          end
          if(_zz_2[2414]) begin
            regVec_2414 <= _zz_regVec_0_1;
          end
          if(_zz_2[2415]) begin
            regVec_2415 <= _zz_regVec_0_1;
          end
          if(_zz_2[2416]) begin
            regVec_2416 <= _zz_regVec_0_1;
          end
          if(_zz_2[2417]) begin
            regVec_2417 <= _zz_regVec_0_1;
          end
          if(_zz_2[2418]) begin
            regVec_2418 <= _zz_regVec_0_1;
          end
          if(_zz_2[2419]) begin
            regVec_2419 <= _zz_regVec_0_1;
          end
          if(_zz_2[2420]) begin
            regVec_2420 <= _zz_regVec_0_1;
          end
          if(_zz_2[2421]) begin
            regVec_2421 <= _zz_regVec_0_1;
          end
          if(_zz_2[2422]) begin
            regVec_2422 <= _zz_regVec_0_1;
          end
          if(_zz_2[2423]) begin
            regVec_2423 <= _zz_regVec_0_1;
          end
          if(_zz_2[2424]) begin
            regVec_2424 <= _zz_regVec_0_1;
          end
          if(_zz_2[2425]) begin
            regVec_2425 <= _zz_regVec_0_1;
          end
          if(_zz_2[2426]) begin
            regVec_2426 <= _zz_regVec_0_1;
          end
          if(_zz_2[2427]) begin
            regVec_2427 <= _zz_regVec_0_1;
          end
          if(_zz_2[2428]) begin
            regVec_2428 <= _zz_regVec_0_1;
          end
          if(_zz_2[2429]) begin
            regVec_2429 <= _zz_regVec_0_1;
          end
          if(_zz_2[2430]) begin
            regVec_2430 <= _zz_regVec_0_1;
          end
          if(_zz_2[2431]) begin
            regVec_2431 <= _zz_regVec_0_1;
          end
          if(_zz_2[2432]) begin
            regVec_2432 <= _zz_regVec_0_1;
          end
          if(_zz_2[2433]) begin
            regVec_2433 <= _zz_regVec_0_1;
          end
          if(_zz_2[2434]) begin
            regVec_2434 <= _zz_regVec_0_1;
          end
          if(_zz_2[2435]) begin
            regVec_2435 <= _zz_regVec_0_1;
          end
          if(_zz_2[2436]) begin
            regVec_2436 <= _zz_regVec_0_1;
          end
          if(_zz_2[2437]) begin
            regVec_2437 <= _zz_regVec_0_1;
          end
          if(_zz_2[2438]) begin
            regVec_2438 <= _zz_regVec_0_1;
          end
          if(_zz_2[2439]) begin
            regVec_2439 <= _zz_regVec_0_1;
          end
          if(_zz_2[2440]) begin
            regVec_2440 <= _zz_regVec_0_1;
          end
          if(_zz_2[2441]) begin
            regVec_2441 <= _zz_regVec_0_1;
          end
          if(_zz_2[2442]) begin
            regVec_2442 <= _zz_regVec_0_1;
          end
          if(_zz_2[2443]) begin
            regVec_2443 <= _zz_regVec_0_1;
          end
          if(_zz_2[2444]) begin
            regVec_2444 <= _zz_regVec_0_1;
          end
          if(_zz_2[2445]) begin
            regVec_2445 <= _zz_regVec_0_1;
          end
          if(_zz_2[2446]) begin
            regVec_2446 <= _zz_regVec_0_1;
          end
          if(_zz_2[2447]) begin
            regVec_2447 <= _zz_regVec_0_1;
          end
          if(_zz_2[2448]) begin
            regVec_2448 <= _zz_regVec_0_1;
          end
          if(_zz_2[2449]) begin
            regVec_2449 <= _zz_regVec_0_1;
          end
          if(_zz_2[2450]) begin
            regVec_2450 <= _zz_regVec_0_1;
          end
          if(_zz_2[2451]) begin
            regVec_2451 <= _zz_regVec_0_1;
          end
          if(_zz_2[2452]) begin
            regVec_2452 <= _zz_regVec_0_1;
          end
          if(_zz_2[2453]) begin
            regVec_2453 <= _zz_regVec_0_1;
          end
          if(_zz_2[2454]) begin
            regVec_2454 <= _zz_regVec_0_1;
          end
          if(_zz_2[2455]) begin
            regVec_2455 <= _zz_regVec_0_1;
          end
          if(_zz_2[2456]) begin
            regVec_2456 <= _zz_regVec_0_1;
          end
          if(_zz_2[2457]) begin
            regVec_2457 <= _zz_regVec_0_1;
          end
          if(_zz_2[2458]) begin
            regVec_2458 <= _zz_regVec_0_1;
          end
          if(_zz_2[2459]) begin
            regVec_2459 <= _zz_regVec_0_1;
          end
          if(_zz_2[2460]) begin
            regVec_2460 <= _zz_regVec_0_1;
          end
          if(_zz_2[2461]) begin
            regVec_2461 <= _zz_regVec_0_1;
          end
          if(_zz_2[2462]) begin
            regVec_2462 <= _zz_regVec_0_1;
          end
          if(_zz_2[2463]) begin
            regVec_2463 <= _zz_regVec_0_1;
          end
          if(_zz_2[2464]) begin
            regVec_2464 <= _zz_regVec_0_1;
          end
          if(_zz_2[2465]) begin
            regVec_2465 <= _zz_regVec_0_1;
          end
          if(_zz_2[2466]) begin
            regVec_2466 <= _zz_regVec_0_1;
          end
          if(_zz_2[2467]) begin
            regVec_2467 <= _zz_regVec_0_1;
          end
          if(_zz_2[2468]) begin
            regVec_2468 <= _zz_regVec_0_1;
          end
          if(_zz_2[2469]) begin
            regVec_2469 <= _zz_regVec_0_1;
          end
          if(_zz_2[2470]) begin
            regVec_2470 <= _zz_regVec_0_1;
          end
          if(_zz_2[2471]) begin
            regVec_2471 <= _zz_regVec_0_1;
          end
          if(_zz_2[2472]) begin
            regVec_2472 <= _zz_regVec_0_1;
          end
          if(_zz_2[2473]) begin
            regVec_2473 <= _zz_regVec_0_1;
          end
          if(_zz_2[2474]) begin
            regVec_2474 <= _zz_regVec_0_1;
          end
          if(_zz_2[2475]) begin
            regVec_2475 <= _zz_regVec_0_1;
          end
          if(_zz_2[2476]) begin
            regVec_2476 <= _zz_regVec_0_1;
          end
          if(_zz_2[2477]) begin
            regVec_2477 <= _zz_regVec_0_1;
          end
          if(_zz_2[2478]) begin
            regVec_2478 <= _zz_regVec_0_1;
          end
          if(_zz_2[2479]) begin
            regVec_2479 <= _zz_regVec_0_1;
          end
          if(_zz_2[2480]) begin
            regVec_2480 <= _zz_regVec_0_1;
          end
          if(_zz_2[2481]) begin
            regVec_2481 <= _zz_regVec_0_1;
          end
          if(_zz_2[2482]) begin
            regVec_2482 <= _zz_regVec_0_1;
          end
          if(_zz_2[2483]) begin
            regVec_2483 <= _zz_regVec_0_1;
          end
          if(_zz_2[2484]) begin
            regVec_2484 <= _zz_regVec_0_1;
          end
          if(_zz_2[2485]) begin
            regVec_2485 <= _zz_regVec_0_1;
          end
          if(_zz_2[2486]) begin
            regVec_2486 <= _zz_regVec_0_1;
          end
          if(_zz_2[2487]) begin
            regVec_2487 <= _zz_regVec_0_1;
          end
          if(_zz_2[2488]) begin
            regVec_2488 <= _zz_regVec_0_1;
          end
          if(_zz_2[2489]) begin
            regVec_2489 <= _zz_regVec_0_1;
          end
          if(_zz_2[2490]) begin
            regVec_2490 <= _zz_regVec_0_1;
          end
          if(_zz_2[2491]) begin
            regVec_2491 <= _zz_regVec_0_1;
          end
          if(_zz_2[2492]) begin
            regVec_2492 <= _zz_regVec_0_1;
          end
          if(_zz_2[2493]) begin
            regVec_2493 <= _zz_regVec_0_1;
          end
          if(_zz_2[2494]) begin
            regVec_2494 <= _zz_regVec_0_1;
          end
          if(_zz_2[2495]) begin
            regVec_2495 <= _zz_regVec_0_1;
          end
          if(_zz_2[2496]) begin
            regVec_2496 <= _zz_regVec_0_1;
          end
          if(_zz_2[2497]) begin
            regVec_2497 <= _zz_regVec_0_1;
          end
          if(_zz_2[2498]) begin
            regVec_2498 <= _zz_regVec_0_1;
          end
          if(_zz_2[2499]) begin
            regVec_2499 <= _zz_regVec_0_1;
          end
          if(_zz_2[2500]) begin
            regVec_2500 <= _zz_regVec_0_1;
          end
          if(_zz_2[2501]) begin
            regVec_2501 <= _zz_regVec_0_1;
          end
          if(_zz_2[2502]) begin
            regVec_2502 <= _zz_regVec_0_1;
          end
          if(_zz_2[2503]) begin
            regVec_2503 <= _zz_regVec_0_1;
          end
          if(_zz_2[2504]) begin
            regVec_2504 <= _zz_regVec_0_1;
          end
          if(_zz_2[2505]) begin
            regVec_2505 <= _zz_regVec_0_1;
          end
          if(_zz_2[2506]) begin
            regVec_2506 <= _zz_regVec_0_1;
          end
          if(_zz_2[2507]) begin
            regVec_2507 <= _zz_regVec_0_1;
          end
          if(_zz_2[2508]) begin
            regVec_2508 <= _zz_regVec_0_1;
          end
          if(_zz_2[2509]) begin
            regVec_2509 <= _zz_regVec_0_1;
          end
          if(_zz_2[2510]) begin
            regVec_2510 <= _zz_regVec_0_1;
          end
          if(_zz_2[2511]) begin
            regVec_2511 <= _zz_regVec_0_1;
          end
          if(_zz_2[2512]) begin
            regVec_2512 <= _zz_regVec_0_1;
          end
          if(_zz_2[2513]) begin
            regVec_2513 <= _zz_regVec_0_1;
          end
          if(_zz_2[2514]) begin
            regVec_2514 <= _zz_regVec_0_1;
          end
          if(_zz_2[2515]) begin
            regVec_2515 <= _zz_regVec_0_1;
          end
          if(_zz_2[2516]) begin
            regVec_2516 <= _zz_regVec_0_1;
          end
          if(_zz_2[2517]) begin
            regVec_2517 <= _zz_regVec_0_1;
          end
          if(_zz_2[2518]) begin
            regVec_2518 <= _zz_regVec_0_1;
          end
          if(_zz_2[2519]) begin
            regVec_2519 <= _zz_regVec_0_1;
          end
          if(_zz_2[2520]) begin
            regVec_2520 <= _zz_regVec_0_1;
          end
          if(_zz_2[2521]) begin
            regVec_2521 <= _zz_regVec_0_1;
          end
          if(_zz_2[2522]) begin
            regVec_2522 <= _zz_regVec_0_1;
          end
          if(_zz_2[2523]) begin
            regVec_2523 <= _zz_regVec_0_1;
          end
          if(_zz_2[2524]) begin
            regVec_2524 <= _zz_regVec_0_1;
          end
          if(_zz_2[2525]) begin
            regVec_2525 <= _zz_regVec_0_1;
          end
          if(_zz_2[2526]) begin
            regVec_2526 <= _zz_regVec_0_1;
          end
          if(_zz_2[2527]) begin
            regVec_2527 <= _zz_regVec_0_1;
          end
          if(_zz_2[2528]) begin
            regVec_2528 <= _zz_regVec_0_1;
          end
          if(_zz_2[2529]) begin
            regVec_2529 <= _zz_regVec_0_1;
          end
          if(_zz_2[2530]) begin
            regVec_2530 <= _zz_regVec_0_1;
          end
          if(_zz_2[2531]) begin
            regVec_2531 <= _zz_regVec_0_1;
          end
          if(_zz_2[2532]) begin
            regVec_2532 <= _zz_regVec_0_1;
          end
          if(_zz_2[2533]) begin
            regVec_2533 <= _zz_regVec_0_1;
          end
          if(_zz_2[2534]) begin
            regVec_2534 <= _zz_regVec_0_1;
          end
          if(_zz_2[2535]) begin
            regVec_2535 <= _zz_regVec_0_1;
          end
          if(_zz_2[2536]) begin
            regVec_2536 <= _zz_regVec_0_1;
          end
          if(_zz_2[2537]) begin
            regVec_2537 <= _zz_regVec_0_1;
          end
          if(_zz_2[2538]) begin
            regVec_2538 <= _zz_regVec_0_1;
          end
          if(_zz_2[2539]) begin
            regVec_2539 <= _zz_regVec_0_1;
          end
          if(_zz_2[2540]) begin
            regVec_2540 <= _zz_regVec_0_1;
          end
          if(_zz_2[2541]) begin
            regVec_2541 <= _zz_regVec_0_1;
          end
          if(_zz_2[2542]) begin
            regVec_2542 <= _zz_regVec_0_1;
          end
          if(_zz_2[2543]) begin
            regVec_2543 <= _zz_regVec_0_1;
          end
          if(_zz_2[2544]) begin
            regVec_2544 <= _zz_regVec_0_1;
          end
          if(_zz_2[2545]) begin
            regVec_2545 <= _zz_regVec_0_1;
          end
          if(_zz_2[2546]) begin
            regVec_2546 <= _zz_regVec_0_1;
          end
          if(_zz_2[2547]) begin
            regVec_2547 <= _zz_regVec_0_1;
          end
          if(_zz_2[2548]) begin
            regVec_2548 <= _zz_regVec_0_1;
          end
          if(_zz_2[2549]) begin
            regVec_2549 <= _zz_regVec_0_1;
          end
          if(_zz_2[2550]) begin
            regVec_2550 <= _zz_regVec_0_1;
          end
          if(_zz_2[2551]) begin
            regVec_2551 <= _zz_regVec_0_1;
          end
          if(_zz_2[2552]) begin
            regVec_2552 <= _zz_regVec_0_1;
          end
          if(_zz_2[2553]) begin
            regVec_2553 <= _zz_regVec_0_1;
          end
          if(_zz_2[2554]) begin
            regVec_2554 <= _zz_regVec_0_1;
          end
          if(_zz_2[2555]) begin
            regVec_2555 <= _zz_regVec_0_1;
          end
          if(_zz_2[2556]) begin
            regVec_2556 <= _zz_regVec_0_1;
          end
          if(_zz_2[2557]) begin
            regVec_2557 <= _zz_regVec_0_1;
          end
          if(_zz_2[2558]) begin
            regVec_2558 <= _zz_regVec_0_1;
          end
          if(_zz_2[2559]) begin
            regVec_2559 <= _zz_regVec_0_1;
          end
          if(_zz_2[2560]) begin
            regVec_2560 <= _zz_regVec_0_1;
          end
          if(_zz_2[2561]) begin
            regVec_2561 <= _zz_regVec_0_1;
          end
          if(_zz_2[2562]) begin
            regVec_2562 <= _zz_regVec_0_1;
          end
          if(_zz_2[2563]) begin
            regVec_2563 <= _zz_regVec_0_1;
          end
          if(_zz_2[2564]) begin
            regVec_2564 <= _zz_regVec_0_1;
          end
          if(_zz_2[2565]) begin
            regVec_2565 <= _zz_regVec_0_1;
          end
          if(_zz_2[2566]) begin
            regVec_2566 <= _zz_regVec_0_1;
          end
          if(_zz_2[2567]) begin
            regVec_2567 <= _zz_regVec_0_1;
          end
          if(_zz_2[2568]) begin
            regVec_2568 <= _zz_regVec_0_1;
          end
          if(_zz_2[2569]) begin
            regVec_2569 <= _zz_regVec_0_1;
          end
          if(_zz_2[2570]) begin
            regVec_2570 <= _zz_regVec_0_1;
          end
          if(_zz_2[2571]) begin
            regVec_2571 <= _zz_regVec_0_1;
          end
          if(_zz_2[2572]) begin
            regVec_2572 <= _zz_regVec_0_1;
          end
          if(_zz_2[2573]) begin
            regVec_2573 <= _zz_regVec_0_1;
          end
          if(_zz_2[2574]) begin
            regVec_2574 <= _zz_regVec_0_1;
          end
          if(_zz_2[2575]) begin
            regVec_2575 <= _zz_regVec_0_1;
          end
          if(_zz_2[2576]) begin
            regVec_2576 <= _zz_regVec_0_1;
          end
          if(_zz_2[2577]) begin
            regVec_2577 <= _zz_regVec_0_1;
          end
          if(_zz_2[2578]) begin
            regVec_2578 <= _zz_regVec_0_1;
          end
          if(_zz_2[2579]) begin
            regVec_2579 <= _zz_regVec_0_1;
          end
          if(_zz_2[2580]) begin
            regVec_2580 <= _zz_regVec_0_1;
          end
          if(_zz_2[2581]) begin
            regVec_2581 <= _zz_regVec_0_1;
          end
          if(_zz_2[2582]) begin
            regVec_2582 <= _zz_regVec_0_1;
          end
          if(_zz_2[2583]) begin
            regVec_2583 <= _zz_regVec_0_1;
          end
          if(_zz_2[2584]) begin
            regVec_2584 <= _zz_regVec_0_1;
          end
          if(_zz_2[2585]) begin
            regVec_2585 <= _zz_regVec_0_1;
          end
          if(_zz_2[2586]) begin
            regVec_2586 <= _zz_regVec_0_1;
          end
          if(_zz_2[2587]) begin
            regVec_2587 <= _zz_regVec_0_1;
          end
          if(_zz_2[2588]) begin
            regVec_2588 <= _zz_regVec_0_1;
          end
          if(_zz_2[2589]) begin
            regVec_2589 <= _zz_regVec_0_1;
          end
          if(_zz_2[2590]) begin
            regVec_2590 <= _zz_regVec_0_1;
          end
          if(_zz_2[2591]) begin
            regVec_2591 <= _zz_regVec_0_1;
          end
          if(_zz_2[2592]) begin
            regVec_2592 <= _zz_regVec_0_1;
          end
          if(_zz_2[2593]) begin
            regVec_2593 <= _zz_regVec_0_1;
          end
          if(_zz_2[2594]) begin
            regVec_2594 <= _zz_regVec_0_1;
          end
          if(_zz_2[2595]) begin
            regVec_2595 <= _zz_regVec_0_1;
          end
          if(_zz_2[2596]) begin
            regVec_2596 <= _zz_regVec_0_1;
          end
          if(_zz_2[2597]) begin
            regVec_2597 <= _zz_regVec_0_1;
          end
          if(_zz_2[2598]) begin
            regVec_2598 <= _zz_regVec_0_1;
          end
          if(_zz_2[2599]) begin
            regVec_2599 <= _zz_regVec_0_1;
          end
          if(_zz_2[2600]) begin
            regVec_2600 <= _zz_regVec_0_1;
          end
          if(_zz_2[2601]) begin
            regVec_2601 <= _zz_regVec_0_1;
          end
          if(_zz_2[2602]) begin
            regVec_2602 <= _zz_regVec_0_1;
          end
          if(_zz_2[2603]) begin
            regVec_2603 <= _zz_regVec_0_1;
          end
          if(_zz_2[2604]) begin
            regVec_2604 <= _zz_regVec_0_1;
          end
          if(_zz_2[2605]) begin
            regVec_2605 <= _zz_regVec_0_1;
          end
          if(_zz_2[2606]) begin
            regVec_2606 <= _zz_regVec_0_1;
          end
          if(_zz_2[2607]) begin
            regVec_2607 <= _zz_regVec_0_1;
          end
          if(_zz_2[2608]) begin
            regVec_2608 <= _zz_regVec_0_1;
          end
          if(_zz_2[2609]) begin
            regVec_2609 <= _zz_regVec_0_1;
          end
          if(_zz_2[2610]) begin
            regVec_2610 <= _zz_regVec_0_1;
          end
          if(_zz_2[2611]) begin
            regVec_2611 <= _zz_regVec_0_1;
          end
          if(_zz_2[2612]) begin
            regVec_2612 <= _zz_regVec_0_1;
          end
          if(_zz_2[2613]) begin
            regVec_2613 <= _zz_regVec_0_1;
          end
          if(_zz_2[2614]) begin
            regVec_2614 <= _zz_regVec_0_1;
          end
          if(_zz_2[2615]) begin
            regVec_2615 <= _zz_regVec_0_1;
          end
          if(_zz_2[2616]) begin
            regVec_2616 <= _zz_regVec_0_1;
          end
          if(_zz_2[2617]) begin
            regVec_2617 <= _zz_regVec_0_1;
          end
          if(_zz_2[2618]) begin
            regVec_2618 <= _zz_regVec_0_1;
          end
          if(_zz_2[2619]) begin
            regVec_2619 <= _zz_regVec_0_1;
          end
          if(_zz_2[2620]) begin
            regVec_2620 <= _zz_regVec_0_1;
          end
          if(_zz_2[2621]) begin
            regVec_2621 <= _zz_regVec_0_1;
          end
          if(_zz_2[2622]) begin
            regVec_2622 <= _zz_regVec_0_1;
          end
          if(_zz_2[2623]) begin
            regVec_2623 <= _zz_regVec_0_1;
          end
          if(_zz_2[2624]) begin
            regVec_2624 <= _zz_regVec_0_1;
          end
          if(_zz_2[2625]) begin
            regVec_2625 <= _zz_regVec_0_1;
          end
          if(_zz_2[2626]) begin
            regVec_2626 <= _zz_regVec_0_1;
          end
          if(_zz_2[2627]) begin
            regVec_2627 <= _zz_regVec_0_1;
          end
          if(_zz_2[2628]) begin
            regVec_2628 <= _zz_regVec_0_1;
          end
          if(_zz_2[2629]) begin
            regVec_2629 <= _zz_regVec_0_1;
          end
          if(_zz_2[2630]) begin
            regVec_2630 <= _zz_regVec_0_1;
          end
          if(_zz_2[2631]) begin
            regVec_2631 <= _zz_regVec_0_1;
          end
          if(_zz_2[2632]) begin
            regVec_2632 <= _zz_regVec_0_1;
          end
          if(_zz_2[2633]) begin
            regVec_2633 <= _zz_regVec_0_1;
          end
          if(_zz_2[2634]) begin
            regVec_2634 <= _zz_regVec_0_1;
          end
          if(_zz_2[2635]) begin
            regVec_2635 <= _zz_regVec_0_1;
          end
          if(_zz_2[2636]) begin
            regVec_2636 <= _zz_regVec_0_1;
          end
          if(_zz_2[2637]) begin
            regVec_2637 <= _zz_regVec_0_1;
          end
          if(_zz_2[2638]) begin
            regVec_2638 <= _zz_regVec_0_1;
          end
          if(_zz_2[2639]) begin
            regVec_2639 <= _zz_regVec_0_1;
          end
          if(_zz_2[2640]) begin
            regVec_2640 <= _zz_regVec_0_1;
          end
          if(_zz_2[2641]) begin
            regVec_2641 <= _zz_regVec_0_1;
          end
          if(_zz_2[2642]) begin
            regVec_2642 <= _zz_regVec_0_1;
          end
          if(_zz_2[2643]) begin
            regVec_2643 <= _zz_regVec_0_1;
          end
          if(_zz_2[2644]) begin
            regVec_2644 <= _zz_regVec_0_1;
          end
          if(_zz_2[2645]) begin
            regVec_2645 <= _zz_regVec_0_1;
          end
          if(_zz_2[2646]) begin
            regVec_2646 <= _zz_regVec_0_1;
          end
          if(_zz_2[2647]) begin
            regVec_2647 <= _zz_regVec_0_1;
          end
          if(_zz_2[2648]) begin
            regVec_2648 <= _zz_regVec_0_1;
          end
          if(_zz_2[2649]) begin
            regVec_2649 <= _zz_regVec_0_1;
          end
          if(_zz_2[2650]) begin
            regVec_2650 <= _zz_regVec_0_1;
          end
          if(_zz_2[2651]) begin
            regVec_2651 <= _zz_regVec_0_1;
          end
          if(_zz_2[2652]) begin
            regVec_2652 <= _zz_regVec_0_1;
          end
          if(_zz_2[2653]) begin
            regVec_2653 <= _zz_regVec_0_1;
          end
          if(_zz_2[2654]) begin
            regVec_2654 <= _zz_regVec_0_1;
          end
          if(_zz_2[2655]) begin
            regVec_2655 <= _zz_regVec_0_1;
          end
          if(_zz_2[2656]) begin
            regVec_2656 <= _zz_regVec_0_1;
          end
          if(_zz_2[2657]) begin
            regVec_2657 <= _zz_regVec_0_1;
          end
          if(_zz_2[2658]) begin
            regVec_2658 <= _zz_regVec_0_1;
          end
          if(_zz_2[2659]) begin
            regVec_2659 <= _zz_regVec_0_1;
          end
          if(_zz_2[2660]) begin
            regVec_2660 <= _zz_regVec_0_1;
          end
          if(_zz_2[2661]) begin
            regVec_2661 <= _zz_regVec_0_1;
          end
          if(_zz_2[2662]) begin
            regVec_2662 <= _zz_regVec_0_1;
          end
          if(_zz_2[2663]) begin
            regVec_2663 <= _zz_regVec_0_1;
          end
          if(_zz_2[2664]) begin
            regVec_2664 <= _zz_regVec_0_1;
          end
          if(_zz_2[2665]) begin
            regVec_2665 <= _zz_regVec_0_1;
          end
          if(_zz_2[2666]) begin
            regVec_2666 <= _zz_regVec_0_1;
          end
          if(_zz_2[2667]) begin
            regVec_2667 <= _zz_regVec_0_1;
          end
          if(_zz_2[2668]) begin
            regVec_2668 <= _zz_regVec_0_1;
          end
          if(_zz_2[2669]) begin
            regVec_2669 <= _zz_regVec_0_1;
          end
          if(_zz_2[2670]) begin
            regVec_2670 <= _zz_regVec_0_1;
          end
          if(_zz_2[2671]) begin
            regVec_2671 <= _zz_regVec_0_1;
          end
          if(_zz_2[2672]) begin
            regVec_2672 <= _zz_regVec_0_1;
          end
          if(_zz_2[2673]) begin
            regVec_2673 <= _zz_regVec_0_1;
          end
          if(_zz_2[2674]) begin
            regVec_2674 <= _zz_regVec_0_1;
          end
          if(_zz_2[2675]) begin
            regVec_2675 <= _zz_regVec_0_1;
          end
          if(_zz_2[2676]) begin
            regVec_2676 <= _zz_regVec_0_1;
          end
          if(_zz_2[2677]) begin
            regVec_2677 <= _zz_regVec_0_1;
          end
          if(_zz_2[2678]) begin
            regVec_2678 <= _zz_regVec_0_1;
          end
          if(_zz_2[2679]) begin
            regVec_2679 <= _zz_regVec_0_1;
          end
          if(_zz_2[2680]) begin
            regVec_2680 <= _zz_regVec_0_1;
          end
          if(_zz_2[2681]) begin
            regVec_2681 <= _zz_regVec_0_1;
          end
          if(_zz_2[2682]) begin
            regVec_2682 <= _zz_regVec_0_1;
          end
          if(_zz_2[2683]) begin
            regVec_2683 <= _zz_regVec_0_1;
          end
          if(_zz_2[2684]) begin
            regVec_2684 <= _zz_regVec_0_1;
          end
          if(_zz_2[2685]) begin
            regVec_2685 <= _zz_regVec_0_1;
          end
          if(_zz_2[2686]) begin
            regVec_2686 <= _zz_regVec_0_1;
          end
          if(_zz_2[2687]) begin
            regVec_2687 <= _zz_regVec_0_1;
          end
          if(_zz_2[2688]) begin
            regVec_2688 <= _zz_regVec_0_1;
          end
          if(_zz_2[2689]) begin
            regVec_2689 <= _zz_regVec_0_1;
          end
          if(_zz_2[2690]) begin
            regVec_2690 <= _zz_regVec_0_1;
          end
          if(_zz_2[2691]) begin
            regVec_2691 <= _zz_regVec_0_1;
          end
          if(_zz_2[2692]) begin
            regVec_2692 <= _zz_regVec_0_1;
          end
          if(_zz_2[2693]) begin
            regVec_2693 <= _zz_regVec_0_1;
          end
          if(_zz_2[2694]) begin
            regVec_2694 <= _zz_regVec_0_1;
          end
          if(_zz_2[2695]) begin
            regVec_2695 <= _zz_regVec_0_1;
          end
          if(_zz_2[2696]) begin
            regVec_2696 <= _zz_regVec_0_1;
          end
          if(_zz_2[2697]) begin
            regVec_2697 <= _zz_regVec_0_1;
          end
          if(_zz_2[2698]) begin
            regVec_2698 <= _zz_regVec_0_1;
          end
          if(_zz_2[2699]) begin
            regVec_2699 <= _zz_regVec_0_1;
          end
          if(_zz_2[2700]) begin
            regVec_2700 <= _zz_regVec_0_1;
          end
          if(_zz_2[2701]) begin
            regVec_2701 <= _zz_regVec_0_1;
          end
          if(_zz_2[2702]) begin
            regVec_2702 <= _zz_regVec_0_1;
          end
          if(_zz_2[2703]) begin
            regVec_2703 <= _zz_regVec_0_1;
          end
          if(_zz_2[2704]) begin
            regVec_2704 <= _zz_regVec_0_1;
          end
          if(_zz_2[2705]) begin
            regVec_2705 <= _zz_regVec_0_1;
          end
          if(_zz_2[2706]) begin
            regVec_2706 <= _zz_regVec_0_1;
          end
          if(_zz_2[2707]) begin
            regVec_2707 <= _zz_regVec_0_1;
          end
          if(_zz_2[2708]) begin
            regVec_2708 <= _zz_regVec_0_1;
          end
          if(_zz_2[2709]) begin
            regVec_2709 <= _zz_regVec_0_1;
          end
          if(_zz_2[2710]) begin
            regVec_2710 <= _zz_regVec_0_1;
          end
          if(_zz_2[2711]) begin
            regVec_2711 <= _zz_regVec_0_1;
          end
          if(_zz_2[2712]) begin
            regVec_2712 <= _zz_regVec_0_1;
          end
          if(_zz_2[2713]) begin
            regVec_2713 <= _zz_regVec_0_1;
          end
          if(_zz_2[2714]) begin
            regVec_2714 <= _zz_regVec_0_1;
          end
          if(_zz_2[2715]) begin
            regVec_2715 <= _zz_regVec_0_1;
          end
          if(_zz_2[2716]) begin
            regVec_2716 <= _zz_regVec_0_1;
          end
          if(_zz_2[2717]) begin
            regVec_2717 <= _zz_regVec_0_1;
          end
          if(_zz_2[2718]) begin
            regVec_2718 <= _zz_regVec_0_1;
          end
          if(_zz_2[2719]) begin
            regVec_2719 <= _zz_regVec_0_1;
          end
          if(_zz_2[2720]) begin
            regVec_2720 <= _zz_regVec_0_1;
          end
          if(_zz_2[2721]) begin
            regVec_2721 <= _zz_regVec_0_1;
          end
          if(_zz_2[2722]) begin
            regVec_2722 <= _zz_regVec_0_1;
          end
          if(_zz_2[2723]) begin
            regVec_2723 <= _zz_regVec_0_1;
          end
          if(_zz_2[2724]) begin
            regVec_2724 <= _zz_regVec_0_1;
          end
          if(_zz_2[2725]) begin
            regVec_2725 <= _zz_regVec_0_1;
          end
          if(_zz_2[2726]) begin
            regVec_2726 <= _zz_regVec_0_1;
          end
          if(_zz_2[2727]) begin
            regVec_2727 <= _zz_regVec_0_1;
          end
          if(_zz_2[2728]) begin
            regVec_2728 <= _zz_regVec_0_1;
          end
          if(_zz_2[2729]) begin
            regVec_2729 <= _zz_regVec_0_1;
          end
          if(_zz_2[2730]) begin
            regVec_2730 <= _zz_regVec_0_1;
          end
          if(_zz_2[2731]) begin
            regVec_2731 <= _zz_regVec_0_1;
          end
          if(_zz_2[2732]) begin
            regVec_2732 <= _zz_regVec_0_1;
          end
          if(_zz_2[2733]) begin
            regVec_2733 <= _zz_regVec_0_1;
          end
          if(_zz_2[2734]) begin
            regVec_2734 <= _zz_regVec_0_1;
          end
          if(_zz_2[2735]) begin
            regVec_2735 <= _zz_regVec_0_1;
          end
          if(_zz_2[2736]) begin
            regVec_2736 <= _zz_regVec_0_1;
          end
          if(_zz_2[2737]) begin
            regVec_2737 <= _zz_regVec_0_1;
          end
          if(_zz_2[2738]) begin
            regVec_2738 <= _zz_regVec_0_1;
          end
          if(_zz_2[2739]) begin
            regVec_2739 <= _zz_regVec_0_1;
          end
          if(_zz_2[2740]) begin
            regVec_2740 <= _zz_regVec_0_1;
          end
          if(_zz_2[2741]) begin
            regVec_2741 <= _zz_regVec_0_1;
          end
          if(_zz_2[2742]) begin
            regVec_2742 <= _zz_regVec_0_1;
          end
          if(_zz_2[2743]) begin
            regVec_2743 <= _zz_regVec_0_1;
          end
          if(_zz_2[2744]) begin
            regVec_2744 <= _zz_regVec_0_1;
          end
          if(_zz_2[2745]) begin
            regVec_2745 <= _zz_regVec_0_1;
          end
          if(_zz_2[2746]) begin
            regVec_2746 <= _zz_regVec_0_1;
          end
          if(_zz_2[2747]) begin
            regVec_2747 <= _zz_regVec_0_1;
          end
          if(_zz_2[2748]) begin
            regVec_2748 <= _zz_regVec_0_1;
          end
          if(_zz_2[2749]) begin
            regVec_2749 <= _zz_regVec_0_1;
          end
          if(_zz_2[2750]) begin
            regVec_2750 <= _zz_regVec_0_1;
          end
          if(_zz_2[2751]) begin
            regVec_2751 <= _zz_regVec_0_1;
          end
          if(_zz_2[2752]) begin
            regVec_2752 <= _zz_regVec_0_1;
          end
          if(_zz_2[2753]) begin
            regVec_2753 <= _zz_regVec_0_1;
          end
          if(_zz_2[2754]) begin
            regVec_2754 <= _zz_regVec_0_1;
          end
          if(_zz_2[2755]) begin
            regVec_2755 <= _zz_regVec_0_1;
          end
          if(_zz_2[2756]) begin
            regVec_2756 <= _zz_regVec_0_1;
          end
          if(_zz_2[2757]) begin
            regVec_2757 <= _zz_regVec_0_1;
          end
          if(_zz_2[2758]) begin
            regVec_2758 <= _zz_regVec_0_1;
          end
          if(_zz_2[2759]) begin
            regVec_2759 <= _zz_regVec_0_1;
          end
          if(_zz_2[2760]) begin
            regVec_2760 <= _zz_regVec_0_1;
          end
          if(_zz_2[2761]) begin
            regVec_2761 <= _zz_regVec_0_1;
          end
          if(_zz_2[2762]) begin
            regVec_2762 <= _zz_regVec_0_1;
          end
          if(_zz_2[2763]) begin
            regVec_2763 <= _zz_regVec_0_1;
          end
          if(_zz_2[2764]) begin
            regVec_2764 <= _zz_regVec_0_1;
          end
          if(_zz_2[2765]) begin
            regVec_2765 <= _zz_regVec_0_1;
          end
          if(_zz_2[2766]) begin
            regVec_2766 <= _zz_regVec_0_1;
          end
          if(_zz_2[2767]) begin
            regVec_2767 <= _zz_regVec_0_1;
          end
          if(_zz_2[2768]) begin
            regVec_2768 <= _zz_regVec_0_1;
          end
          if(_zz_2[2769]) begin
            regVec_2769 <= _zz_regVec_0_1;
          end
          if(_zz_2[2770]) begin
            regVec_2770 <= _zz_regVec_0_1;
          end
          if(_zz_2[2771]) begin
            regVec_2771 <= _zz_regVec_0_1;
          end
          if(_zz_2[2772]) begin
            regVec_2772 <= _zz_regVec_0_1;
          end
          if(_zz_2[2773]) begin
            regVec_2773 <= _zz_regVec_0_1;
          end
          if(_zz_2[2774]) begin
            regVec_2774 <= _zz_regVec_0_1;
          end
          if(_zz_2[2775]) begin
            regVec_2775 <= _zz_regVec_0_1;
          end
          if(_zz_2[2776]) begin
            regVec_2776 <= _zz_regVec_0_1;
          end
          if(_zz_2[2777]) begin
            regVec_2777 <= _zz_regVec_0_1;
          end
          if(_zz_2[2778]) begin
            regVec_2778 <= _zz_regVec_0_1;
          end
          if(_zz_2[2779]) begin
            regVec_2779 <= _zz_regVec_0_1;
          end
          if(_zz_2[2780]) begin
            regVec_2780 <= _zz_regVec_0_1;
          end
          if(_zz_2[2781]) begin
            regVec_2781 <= _zz_regVec_0_1;
          end
          if(_zz_2[2782]) begin
            regVec_2782 <= _zz_regVec_0_1;
          end
          if(_zz_2[2783]) begin
            regVec_2783 <= _zz_regVec_0_1;
          end
          if(_zz_2[2784]) begin
            regVec_2784 <= _zz_regVec_0_1;
          end
          if(_zz_2[2785]) begin
            regVec_2785 <= _zz_regVec_0_1;
          end
          if(_zz_2[2786]) begin
            regVec_2786 <= _zz_regVec_0_1;
          end
          if(_zz_2[2787]) begin
            regVec_2787 <= _zz_regVec_0_1;
          end
          if(_zz_2[2788]) begin
            regVec_2788 <= _zz_regVec_0_1;
          end
          if(_zz_2[2789]) begin
            regVec_2789 <= _zz_regVec_0_1;
          end
          if(_zz_2[2790]) begin
            regVec_2790 <= _zz_regVec_0_1;
          end
          if(_zz_2[2791]) begin
            regVec_2791 <= _zz_regVec_0_1;
          end
          if(_zz_2[2792]) begin
            regVec_2792 <= _zz_regVec_0_1;
          end
          if(_zz_2[2793]) begin
            regVec_2793 <= _zz_regVec_0_1;
          end
          if(_zz_2[2794]) begin
            regVec_2794 <= _zz_regVec_0_1;
          end
          if(_zz_2[2795]) begin
            regVec_2795 <= _zz_regVec_0_1;
          end
          if(_zz_2[2796]) begin
            regVec_2796 <= _zz_regVec_0_1;
          end
          if(_zz_2[2797]) begin
            regVec_2797 <= _zz_regVec_0_1;
          end
          if(_zz_2[2798]) begin
            regVec_2798 <= _zz_regVec_0_1;
          end
          if(_zz_2[2799]) begin
            regVec_2799 <= _zz_regVec_0_1;
          end
          if(_zz_2[2800]) begin
            regVec_2800 <= _zz_regVec_0_1;
          end
          if(_zz_2[2801]) begin
            regVec_2801 <= _zz_regVec_0_1;
          end
          if(_zz_2[2802]) begin
            regVec_2802 <= _zz_regVec_0_1;
          end
          if(_zz_2[2803]) begin
            regVec_2803 <= _zz_regVec_0_1;
          end
          if(_zz_2[2804]) begin
            regVec_2804 <= _zz_regVec_0_1;
          end
          if(_zz_2[2805]) begin
            regVec_2805 <= _zz_regVec_0_1;
          end
          if(_zz_2[2806]) begin
            regVec_2806 <= _zz_regVec_0_1;
          end
          if(_zz_2[2807]) begin
            regVec_2807 <= _zz_regVec_0_1;
          end
          if(_zz_2[2808]) begin
            regVec_2808 <= _zz_regVec_0_1;
          end
          if(_zz_2[2809]) begin
            regVec_2809 <= _zz_regVec_0_1;
          end
          if(_zz_2[2810]) begin
            regVec_2810 <= _zz_regVec_0_1;
          end
          if(_zz_2[2811]) begin
            regVec_2811 <= _zz_regVec_0_1;
          end
          if(_zz_2[2812]) begin
            regVec_2812 <= _zz_regVec_0_1;
          end
          if(_zz_2[2813]) begin
            regVec_2813 <= _zz_regVec_0_1;
          end
          if(_zz_2[2814]) begin
            regVec_2814 <= _zz_regVec_0_1;
          end
          if(_zz_2[2815]) begin
            regVec_2815 <= _zz_regVec_0_1;
          end
          if(_zz_2[2816]) begin
            regVec_2816 <= _zz_regVec_0_1;
          end
          if(_zz_2[2817]) begin
            regVec_2817 <= _zz_regVec_0_1;
          end
          if(_zz_2[2818]) begin
            regVec_2818 <= _zz_regVec_0_1;
          end
          if(_zz_2[2819]) begin
            regVec_2819 <= _zz_regVec_0_1;
          end
          if(_zz_2[2820]) begin
            regVec_2820 <= _zz_regVec_0_1;
          end
          if(_zz_2[2821]) begin
            regVec_2821 <= _zz_regVec_0_1;
          end
          if(_zz_2[2822]) begin
            regVec_2822 <= _zz_regVec_0_1;
          end
          if(_zz_2[2823]) begin
            regVec_2823 <= _zz_regVec_0_1;
          end
          if(_zz_2[2824]) begin
            regVec_2824 <= _zz_regVec_0_1;
          end
          if(_zz_2[2825]) begin
            regVec_2825 <= _zz_regVec_0_1;
          end
          if(_zz_2[2826]) begin
            regVec_2826 <= _zz_regVec_0_1;
          end
          if(_zz_2[2827]) begin
            regVec_2827 <= _zz_regVec_0_1;
          end
          if(_zz_2[2828]) begin
            regVec_2828 <= _zz_regVec_0_1;
          end
          if(_zz_2[2829]) begin
            regVec_2829 <= _zz_regVec_0_1;
          end
          if(_zz_2[2830]) begin
            regVec_2830 <= _zz_regVec_0_1;
          end
          if(_zz_2[2831]) begin
            regVec_2831 <= _zz_regVec_0_1;
          end
          if(_zz_2[2832]) begin
            regVec_2832 <= _zz_regVec_0_1;
          end
          if(_zz_2[2833]) begin
            regVec_2833 <= _zz_regVec_0_1;
          end
          if(_zz_2[2834]) begin
            regVec_2834 <= _zz_regVec_0_1;
          end
          if(_zz_2[2835]) begin
            regVec_2835 <= _zz_regVec_0_1;
          end
          if(_zz_2[2836]) begin
            regVec_2836 <= _zz_regVec_0_1;
          end
          if(_zz_2[2837]) begin
            regVec_2837 <= _zz_regVec_0_1;
          end
          if(_zz_2[2838]) begin
            regVec_2838 <= _zz_regVec_0_1;
          end
          if(_zz_2[2839]) begin
            regVec_2839 <= _zz_regVec_0_1;
          end
          if(_zz_2[2840]) begin
            regVec_2840 <= _zz_regVec_0_1;
          end
          if(_zz_2[2841]) begin
            regVec_2841 <= _zz_regVec_0_1;
          end
          if(_zz_2[2842]) begin
            regVec_2842 <= _zz_regVec_0_1;
          end
          if(_zz_2[2843]) begin
            regVec_2843 <= _zz_regVec_0_1;
          end
          if(_zz_2[2844]) begin
            regVec_2844 <= _zz_regVec_0_1;
          end
          if(_zz_2[2845]) begin
            regVec_2845 <= _zz_regVec_0_1;
          end
          if(_zz_2[2846]) begin
            regVec_2846 <= _zz_regVec_0_1;
          end
          if(_zz_2[2847]) begin
            regVec_2847 <= _zz_regVec_0_1;
          end
          if(_zz_2[2848]) begin
            regVec_2848 <= _zz_regVec_0_1;
          end
          if(_zz_2[2849]) begin
            regVec_2849 <= _zz_regVec_0_1;
          end
          if(_zz_2[2850]) begin
            regVec_2850 <= _zz_regVec_0_1;
          end
          if(_zz_2[2851]) begin
            regVec_2851 <= _zz_regVec_0_1;
          end
          if(_zz_2[2852]) begin
            regVec_2852 <= _zz_regVec_0_1;
          end
          if(_zz_2[2853]) begin
            regVec_2853 <= _zz_regVec_0_1;
          end
          if(_zz_2[2854]) begin
            regVec_2854 <= _zz_regVec_0_1;
          end
          if(_zz_2[2855]) begin
            regVec_2855 <= _zz_regVec_0_1;
          end
          if(_zz_2[2856]) begin
            regVec_2856 <= _zz_regVec_0_1;
          end
          if(_zz_2[2857]) begin
            regVec_2857 <= _zz_regVec_0_1;
          end
          if(_zz_2[2858]) begin
            regVec_2858 <= _zz_regVec_0_1;
          end
          if(_zz_2[2859]) begin
            regVec_2859 <= _zz_regVec_0_1;
          end
          if(_zz_2[2860]) begin
            regVec_2860 <= _zz_regVec_0_1;
          end
          if(_zz_2[2861]) begin
            regVec_2861 <= _zz_regVec_0_1;
          end
          if(_zz_2[2862]) begin
            regVec_2862 <= _zz_regVec_0_1;
          end
          if(_zz_2[2863]) begin
            regVec_2863 <= _zz_regVec_0_1;
          end
          if(_zz_2[2864]) begin
            regVec_2864 <= _zz_regVec_0_1;
          end
          if(_zz_2[2865]) begin
            regVec_2865 <= _zz_regVec_0_1;
          end
          if(_zz_2[2866]) begin
            regVec_2866 <= _zz_regVec_0_1;
          end
          if(_zz_2[2867]) begin
            regVec_2867 <= _zz_regVec_0_1;
          end
          if(_zz_2[2868]) begin
            regVec_2868 <= _zz_regVec_0_1;
          end
          if(_zz_2[2869]) begin
            regVec_2869 <= _zz_regVec_0_1;
          end
          if(_zz_2[2870]) begin
            regVec_2870 <= _zz_regVec_0_1;
          end
          if(_zz_2[2871]) begin
            regVec_2871 <= _zz_regVec_0_1;
          end
          if(_zz_2[2872]) begin
            regVec_2872 <= _zz_regVec_0_1;
          end
          if(_zz_2[2873]) begin
            regVec_2873 <= _zz_regVec_0_1;
          end
          if(_zz_2[2874]) begin
            regVec_2874 <= _zz_regVec_0_1;
          end
          if(_zz_2[2875]) begin
            regVec_2875 <= _zz_regVec_0_1;
          end
          if(_zz_2[2876]) begin
            regVec_2876 <= _zz_regVec_0_1;
          end
          if(_zz_2[2877]) begin
            regVec_2877 <= _zz_regVec_0_1;
          end
          if(_zz_2[2878]) begin
            regVec_2878 <= _zz_regVec_0_1;
          end
          if(_zz_2[2879]) begin
            regVec_2879 <= _zz_regVec_0_1;
          end
          if(_zz_2[2880]) begin
            regVec_2880 <= _zz_regVec_0_1;
          end
          if(_zz_2[2881]) begin
            regVec_2881 <= _zz_regVec_0_1;
          end
          if(_zz_2[2882]) begin
            regVec_2882 <= _zz_regVec_0_1;
          end
          if(_zz_2[2883]) begin
            regVec_2883 <= _zz_regVec_0_1;
          end
          if(_zz_2[2884]) begin
            regVec_2884 <= _zz_regVec_0_1;
          end
          if(_zz_2[2885]) begin
            regVec_2885 <= _zz_regVec_0_1;
          end
          if(_zz_2[2886]) begin
            regVec_2886 <= _zz_regVec_0_1;
          end
          if(_zz_2[2887]) begin
            regVec_2887 <= _zz_regVec_0_1;
          end
          if(_zz_2[2888]) begin
            regVec_2888 <= _zz_regVec_0_1;
          end
          if(_zz_2[2889]) begin
            regVec_2889 <= _zz_regVec_0_1;
          end
          if(_zz_2[2890]) begin
            regVec_2890 <= _zz_regVec_0_1;
          end
          if(_zz_2[2891]) begin
            regVec_2891 <= _zz_regVec_0_1;
          end
          if(_zz_2[2892]) begin
            regVec_2892 <= _zz_regVec_0_1;
          end
          if(_zz_2[2893]) begin
            regVec_2893 <= _zz_regVec_0_1;
          end
          if(_zz_2[2894]) begin
            regVec_2894 <= _zz_regVec_0_1;
          end
          if(_zz_2[2895]) begin
            regVec_2895 <= _zz_regVec_0_1;
          end
          if(_zz_2[2896]) begin
            regVec_2896 <= _zz_regVec_0_1;
          end
          if(_zz_2[2897]) begin
            regVec_2897 <= _zz_regVec_0_1;
          end
          if(_zz_2[2898]) begin
            regVec_2898 <= _zz_regVec_0_1;
          end
          if(_zz_2[2899]) begin
            regVec_2899 <= _zz_regVec_0_1;
          end
          if(_zz_2[2900]) begin
            regVec_2900 <= _zz_regVec_0_1;
          end
          if(_zz_2[2901]) begin
            regVec_2901 <= _zz_regVec_0_1;
          end
          if(_zz_2[2902]) begin
            regVec_2902 <= _zz_regVec_0_1;
          end
          if(_zz_2[2903]) begin
            regVec_2903 <= _zz_regVec_0_1;
          end
          if(_zz_2[2904]) begin
            regVec_2904 <= _zz_regVec_0_1;
          end
          if(_zz_2[2905]) begin
            regVec_2905 <= _zz_regVec_0_1;
          end
          if(_zz_2[2906]) begin
            regVec_2906 <= _zz_regVec_0_1;
          end
          if(_zz_2[2907]) begin
            regVec_2907 <= _zz_regVec_0_1;
          end
          if(_zz_2[2908]) begin
            regVec_2908 <= _zz_regVec_0_1;
          end
          if(_zz_2[2909]) begin
            regVec_2909 <= _zz_regVec_0_1;
          end
          if(_zz_2[2910]) begin
            regVec_2910 <= _zz_regVec_0_1;
          end
          if(_zz_2[2911]) begin
            regVec_2911 <= _zz_regVec_0_1;
          end
          if(_zz_2[2912]) begin
            regVec_2912 <= _zz_regVec_0_1;
          end
          if(_zz_2[2913]) begin
            regVec_2913 <= _zz_regVec_0_1;
          end
          if(_zz_2[2914]) begin
            regVec_2914 <= _zz_regVec_0_1;
          end
          if(_zz_2[2915]) begin
            regVec_2915 <= _zz_regVec_0_1;
          end
          if(_zz_2[2916]) begin
            regVec_2916 <= _zz_regVec_0_1;
          end
          if(_zz_2[2917]) begin
            regVec_2917 <= _zz_regVec_0_1;
          end
          if(_zz_2[2918]) begin
            regVec_2918 <= _zz_regVec_0_1;
          end
          if(_zz_2[2919]) begin
            regVec_2919 <= _zz_regVec_0_1;
          end
          if(_zz_2[2920]) begin
            regVec_2920 <= _zz_regVec_0_1;
          end
          if(_zz_2[2921]) begin
            regVec_2921 <= _zz_regVec_0_1;
          end
          if(_zz_2[2922]) begin
            regVec_2922 <= _zz_regVec_0_1;
          end
          if(_zz_2[2923]) begin
            regVec_2923 <= _zz_regVec_0_1;
          end
          if(_zz_2[2924]) begin
            regVec_2924 <= _zz_regVec_0_1;
          end
          if(_zz_2[2925]) begin
            regVec_2925 <= _zz_regVec_0_1;
          end
          if(_zz_2[2926]) begin
            regVec_2926 <= _zz_regVec_0_1;
          end
          if(_zz_2[2927]) begin
            regVec_2927 <= _zz_regVec_0_1;
          end
          if(_zz_2[2928]) begin
            regVec_2928 <= _zz_regVec_0_1;
          end
          if(_zz_2[2929]) begin
            regVec_2929 <= _zz_regVec_0_1;
          end
          if(_zz_2[2930]) begin
            regVec_2930 <= _zz_regVec_0_1;
          end
          if(_zz_2[2931]) begin
            regVec_2931 <= _zz_regVec_0_1;
          end
          if(_zz_2[2932]) begin
            regVec_2932 <= _zz_regVec_0_1;
          end
          if(_zz_2[2933]) begin
            regVec_2933 <= _zz_regVec_0_1;
          end
          if(_zz_2[2934]) begin
            regVec_2934 <= _zz_regVec_0_1;
          end
          if(_zz_2[2935]) begin
            regVec_2935 <= _zz_regVec_0_1;
          end
          if(_zz_2[2936]) begin
            regVec_2936 <= _zz_regVec_0_1;
          end
          if(_zz_2[2937]) begin
            regVec_2937 <= _zz_regVec_0_1;
          end
          if(_zz_2[2938]) begin
            regVec_2938 <= _zz_regVec_0_1;
          end
          if(_zz_2[2939]) begin
            regVec_2939 <= _zz_regVec_0_1;
          end
          if(_zz_2[2940]) begin
            regVec_2940 <= _zz_regVec_0_1;
          end
          if(_zz_2[2941]) begin
            regVec_2941 <= _zz_regVec_0_1;
          end
          if(_zz_2[2942]) begin
            regVec_2942 <= _zz_regVec_0_1;
          end
          if(_zz_2[2943]) begin
            regVec_2943 <= _zz_regVec_0_1;
          end
          if(_zz_2[2944]) begin
            regVec_2944 <= _zz_regVec_0_1;
          end
          if(_zz_2[2945]) begin
            regVec_2945 <= _zz_regVec_0_1;
          end
          if(_zz_2[2946]) begin
            regVec_2946 <= _zz_regVec_0_1;
          end
          if(_zz_2[2947]) begin
            regVec_2947 <= _zz_regVec_0_1;
          end
          if(_zz_2[2948]) begin
            regVec_2948 <= _zz_regVec_0_1;
          end
          if(_zz_2[2949]) begin
            regVec_2949 <= _zz_regVec_0_1;
          end
          if(_zz_2[2950]) begin
            regVec_2950 <= _zz_regVec_0_1;
          end
          if(_zz_2[2951]) begin
            regVec_2951 <= _zz_regVec_0_1;
          end
          if(_zz_2[2952]) begin
            regVec_2952 <= _zz_regVec_0_1;
          end
          if(_zz_2[2953]) begin
            regVec_2953 <= _zz_regVec_0_1;
          end
          if(_zz_2[2954]) begin
            regVec_2954 <= _zz_regVec_0_1;
          end
          if(_zz_2[2955]) begin
            regVec_2955 <= _zz_regVec_0_1;
          end
          if(_zz_2[2956]) begin
            regVec_2956 <= _zz_regVec_0_1;
          end
          if(_zz_2[2957]) begin
            regVec_2957 <= _zz_regVec_0_1;
          end
          if(_zz_2[2958]) begin
            regVec_2958 <= _zz_regVec_0_1;
          end
          if(_zz_2[2959]) begin
            regVec_2959 <= _zz_regVec_0_1;
          end
          if(_zz_2[2960]) begin
            regVec_2960 <= _zz_regVec_0_1;
          end
          if(_zz_2[2961]) begin
            regVec_2961 <= _zz_regVec_0_1;
          end
          if(_zz_2[2962]) begin
            regVec_2962 <= _zz_regVec_0_1;
          end
          if(_zz_2[2963]) begin
            regVec_2963 <= _zz_regVec_0_1;
          end
          if(_zz_2[2964]) begin
            regVec_2964 <= _zz_regVec_0_1;
          end
          if(_zz_2[2965]) begin
            regVec_2965 <= _zz_regVec_0_1;
          end
          if(_zz_2[2966]) begin
            regVec_2966 <= _zz_regVec_0_1;
          end
          if(_zz_2[2967]) begin
            regVec_2967 <= _zz_regVec_0_1;
          end
          if(_zz_2[2968]) begin
            regVec_2968 <= _zz_regVec_0_1;
          end
          if(_zz_2[2969]) begin
            regVec_2969 <= _zz_regVec_0_1;
          end
          if(_zz_2[2970]) begin
            regVec_2970 <= _zz_regVec_0_1;
          end
          if(_zz_2[2971]) begin
            regVec_2971 <= _zz_regVec_0_1;
          end
          if(_zz_2[2972]) begin
            regVec_2972 <= _zz_regVec_0_1;
          end
          if(_zz_2[2973]) begin
            regVec_2973 <= _zz_regVec_0_1;
          end
          if(_zz_2[2974]) begin
            regVec_2974 <= _zz_regVec_0_1;
          end
          if(_zz_2[2975]) begin
            regVec_2975 <= _zz_regVec_0_1;
          end
          if(_zz_2[2976]) begin
            regVec_2976 <= _zz_regVec_0_1;
          end
          if(_zz_2[2977]) begin
            regVec_2977 <= _zz_regVec_0_1;
          end
          if(_zz_2[2978]) begin
            regVec_2978 <= _zz_regVec_0_1;
          end
          if(_zz_2[2979]) begin
            regVec_2979 <= _zz_regVec_0_1;
          end
          if(_zz_2[2980]) begin
            regVec_2980 <= _zz_regVec_0_1;
          end
          if(_zz_2[2981]) begin
            regVec_2981 <= _zz_regVec_0_1;
          end
          if(_zz_2[2982]) begin
            regVec_2982 <= _zz_regVec_0_1;
          end
          if(_zz_2[2983]) begin
            regVec_2983 <= _zz_regVec_0_1;
          end
          if(_zz_2[2984]) begin
            regVec_2984 <= _zz_regVec_0_1;
          end
          if(_zz_2[2985]) begin
            regVec_2985 <= _zz_regVec_0_1;
          end
          if(_zz_2[2986]) begin
            regVec_2986 <= _zz_regVec_0_1;
          end
          if(_zz_2[2987]) begin
            regVec_2987 <= _zz_regVec_0_1;
          end
          if(_zz_2[2988]) begin
            regVec_2988 <= _zz_regVec_0_1;
          end
          if(_zz_2[2989]) begin
            regVec_2989 <= _zz_regVec_0_1;
          end
          if(_zz_2[2990]) begin
            regVec_2990 <= _zz_regVec_0_1;
          end
          if(_zz_2[2991]) begin
            regVec_2991 <= _zz_regVec_0_1;
          end
          if(_zz_2[2992]) begin
            regVec_2992 <= _zz_regVec_0_1;
          end
          if(_zz_2[2993]) begin
            regVec_2993 <= _zz_regVec_0_1;
          end
          if(_zz_2[2994]) begin
            regVec_2994 <= _zz_regVec_0_1;
          end
          if(_zz_2[2995]) begin
            regVec_2995 <= _zz_regVec_0_1;
          end
          if(_zz_2[2996]) begin
            regVec_2996 <= _zz_regVec_0_1;
          end
          if(_zz_2[2997]) begin
            regVec_2997 <= _zz_regVec_0_1;
          end
          if(_zz_2[2998]) begin
            regVec_2998 <= _zz_regVec_0_1;
          end
          if(_zz_2[2999]) begin
            regVec_2999 <= _zz_regVec_0_1;
          end
          if(_zz_2[3000]) begin
            regVec_3000 <= _zz_regVec_0_1;
          end
          if(_zz_2[3001]) begin
            regVec_3001 <= _zz_regVec_0_1;
          end
          if(_zz_2[3002]) begin
            regVec_3002 <= _zz_regVec_0_1;
          end
          if(_zz_2[3003]) begin
            regVec_3003 <= _zz_regVec_0_1;
          end
          if(_zz_2[3004]) begin
            regVec_3004 <= _zz_regVec_0_1;
          end
          if(_zz_2[3005]) begin
            regVec_3005 <= _zz_regVec_0_1;
          end
          if(_zz_2[3006]) begin
            regVec_3006 <= _zz_regVec_0_1;
          end
          if(_zz_2[3007]) begin
            regVec_3007 <= _zz_regVec_0_1;
          end
          if(_zz_2[3008]) begin
            regVec_3008 <= _zz_regVec_0_1;
          end
          if(_zz_2[3009]) begin
            regVec_3009 <= _zz_regVec_0_1;
          end
          if(_zz_2[3010]) begin
            regVec_3010 <= _zz_regVec_0_1;
          end
          if(_zz_2[3011]) begin
            regVec_3011 <= _zz_regVec_0_1;
          end
          if(_zz_2[3012]) begin
            regVec_3012 <= _zz_regVec_0_1;
          end
          if(_zz_2[3013]) begin
            regVec_3013 <= _zz_regVec_0_1;
          end
          if(_zz_2[3014]) begin
            regVec_3014 <= _zz_regVec_0_1;
          end
          if(_zz_2[3015]) begin
            regVec_3015 <= _zz_regVec_0_1;
          end
          if(_zz_2[3016]) begin
            regVec_3016 <= _zz_regVec_0_1;
          end
          if(_zz_2[3017]) begin
            regVec_3017 <= _zz_regVec_0_1;
          end
          if(_zz_2[3018]) begin
            regVec_3018 <= _zz_regVec_0_1;
          end
          if(_zz_2[3019]) begin
            regVec_3019 <= _zz_regVec_0_1;
          end
          if(_zz_2[3020]) begin
            regVec_3020 <= _zz_regVec_0_1;
          end
          if(_zz_2[3021]) begin
            regVec_3021 <= _zz_regVec_0_1;
          end
          if(_zz_2[3022]) begin
            regVec_3022 <= _zz_regVec_0_1;
          end
          if(_zz_2[3023]) begin
            regVec_3023 <= _zz_regVec_0_1;
          end
          if(_zz_2[3024]) begin
            regVec_3024 <= _zz_regVec_0_1;
          end
          if(_zz_2[3025]) begin
            regVec_3025 <= _zz_regVec_0_1;
          end
          if(_zz_2[3026]) begin
            regVec_3026 <= _zz_regVec_0_1;
          end
          if(_zz_2[3027]) begin
            regVec_3027 <= _zz_regVec_0_1;
          end
          if(_zz_2[3028]) begin
            regVec_3028 <= _zz_regVec_0_1;
          end
          if(_zz_2[3029]) begin
            regVec_3029 <= _zz_regVec_0_1;
          end
          if(_zz_2[3030]) begin
            regVec_3030 <= _zz_regVec_0_1;
          end
          if(_zz_2[3031]) begin
            regVec_3031 <= _zz_regVec_0_1;
          end
          if(_zz_2[3032]) begin
            regVec_3032 <= _zz_regVec_0_1;
          end
          if(_zz_2[3033]) begin
            regVec_3033 <= _zz_regVec_0_1;
          end
          if(_zz_2[3034]) begin
            regVec_3034 <= _zz_regVec_0_1;
          end
          if(_zz_2[3035]) begin
            regVec_3035 <= _zz_regVec_0_1;
          end
          if(_zz_2[3036]) begin
            regVec_3036 <= _zz_regVec_0_1;
          end
          if(_zz_2[3037]) begin
            regVec_3037 <= _zz_regVec_0_1;
          end
          if(_zz_2[3038]) begin
            regVec_3038 <= _zz_regVec_0_1;
          end
          if(_zz_2[3039]) begin
            regVec_3039 <= _zz_regVec_0_1;
          end
          if(_zz_2[3040]) begin
            regVec_3040 <= _zz_regVec_0_1;
          end
          if(_zz_2[3041]) begin
            regVec_3041 <= _zz_regVec_0_1;
          end
          if(_zz_2[3042]) begin
            regVec_3042 <= _zz_regVec_0_1;
          end
          if(_zz_2[3043]) begin
            regVec_3043 <= _zz_regVec_0_1;
          end
          if(_zz_2[3044]) begin
            regVec_3044 <= _zz_regVec_0_1;
          end
          if(_zz_2[3045]) begin
            regVec_3045 <= _zz_regVec_0_1;
          end
          if(_zz_2[3046]) begin
            regVec_3046 <= _zz_regVec_0_1;
          end
          if(_zz_2[3047]) begin
            regVec_3047 <= _zz_regVec_0_1;
          end
          if(_zz_2[3048]) begin
            regVec_3048 <= _zz_regVec_0_1;
          end
          if(_zz_2[3049]) begin
            regVec_3049 <= _zz_regVec_0_1;
          end
          if(_zz_2[3050]) begin
            regVec_3050 <= _zz_regVec_0_1;
          end
          if(_zz_2[3051]) begin
            regVec_3051 <= _zz_regVec_0_1;
          end
          if(_zz_2[3052]) begin
            regVec_3052 <= _zz_regVec_0_1;
          end
          if(_zz_2[3053]) begin
            regVec_3053 <= _zz_regVec_0_1;
          end
          if(_zz_2[3054]) begin
            regVec_3054 <= _zz_regVec_0_1;
          end
          if(_zz_2[3055]) begin
            regVec_3055 <= _zz_regVec_0_1;
          end
          if(_zz_2[3056]) begin
            regVec_3056 <= _zz_regVec_0_1;
          end
          if(_zz_2[3057]) begin
            regVec_3057 <= _zz_regVec_0_1;
          end
          if(_zz_2[3058]) begin
            regVec_3058 <= _zz_regVec_0_1;
          end
          if(_zz_2[3059]) begin
            regVec_3059 <= _zz_regVec_0_1;
          end
          if(_zz_2[3060]) begin
            regVec_3060 <= _zz_regVec_0_1;
          end
          if(_zz_2[3061]) begin
            regVec_3061 <= _zz_regVec_0_1;
          end
          if(_zz_2[3062]) begin
            regVec_3062 <= _zz_regVec_0_1;
          end
          if(_zz_2[3063]) begin
            regVec_3063 <= _zz_regVec_0_1;
          end
          if(_zz_2[3064]) begin
            regVec_3064 <= _zz_regVec_0_1;
          end
          if(_zz_2[3065]) begin
            regVec_3065 <= _zz_regVec_0_1;
          end
          if(_zz_2[3066]) begin
            regVec_3066 <= _zz_regVec_0_1;
          end
          if(_zz_2[3067]) begin
            regVec_3067 <= _zz_regVec_0_1;
          end
          if(_zz_2[3068]) begin
            regVec_3068 <= _zz_regVec_0_1;
          end
          if(_zz_2[3069]) begin
            regVec_3069 <= _zz_regVec_0_1;
          end
          if(_zz_2[3070]) begin
            regVec_3070 <= _zz_regVec_0_1;
          end
          if(_zz_2[3071]) begin
            regVec_3071 <= _zz_regVec_0_1;
          end
          if(_zz_2[3072]) begin
            regVec_3072 <= _zz_regVec_0_1;
          end
          if(_zz_2[3073]) begin
            regVec_3073 <= _zz_regVec_0_1;
          end
          if(_zz_2[3074]) begin
            regVec_3074 <= _zz_regVec_0_1;
          end
          if(_zz_2[3075]) begin
            regVec_3075 <= _zz_regVec_0_1;
          end
          if(_zz_2[3076]) begin
            regVec_3076 <= _zz_regVec_0_1;
          end
          if(_zz_2[3077]) begin
            regVec_3077 <= _zz_regVec_0_1;
          end
          if(_zz_2[3078]) begin
            regVec_3078 <= _zz_regVec_0_1;
          end
          if(_zz_2[3079]) begin
            regVec_3079 <= _zz_regVec_0_1;
          end
          if(_zz_2[3080]) begin
            regVec_3080 <= _zz_regVec_0_1;
          end
          if(_zz_2[3081]) begin
            regVec_3081 <= _zz_regVec_0_1;
          end
          if(_zz_2[3082]) begin
            regVec_3082 <= _zz_regVec_0_1;
          end
          if(_zz_2[3083]) begin
            regVec_3083 <= _zz_regVec_0_1;
          end
          if(_zz_2[3084]) begin
            regVec_3084 <= _zz_regVec_0_1;
          end
          if(_zz_2[3085]) begin
            regVec_3085 <= _zz_regVec_0_1;
          end
          if(_zz_2[3086]) begin
            regVec_3086 <= _zz_regVec_0_1;
          end
          if(_zz_2[3087]) begin
            regVec_3087 <= _zz_regVec_0_1;
          end
          if(_zz_2[3088]) begin
            regVec_3088 <= _zz_regVec_0_1;
          end
          if(_zz_2[3089]) begin
            regVec_3089 <= _zz_regVec_0_1;
          end
          if(_zz_2[3090]) begin
            regVec_3090 <= _zz_regVec_0_1;
          end
          if(_zz_2[3091]) begin
            regVec_3091 <= _zz_regVec_0_1;
          end
          if(_zz_2[3092]) begin
            regVec_3092 <= _zz_regVec_0_1;
          end
          if(_zz_2[3093]) begin
            regVec_3093 <= _zz_regVec_0_1;
          end
          if(_zz_2[3094]) begin
            regVec_3094 <= _zz_regVec_0_1;
          end
          if(_zz_2[3095]) begin
            regVec_3095 <= _zz_regVec_0_1;
          end
          if(_zz_2[3096]) begin
            regVec_3096 <= _zz_regVec_0_1;
          end
          if(_zz_2[3097]) begin
            regVec_3097 <= _zz_regVec_0_1;
          end
          if(_zz_2[3098]) begin
            regVec_3098 <= _zz_regVec_0_1;
          end
          if(_zz_2[3099]) begin
            regVec_3099 <= _zz_regVec_0_1;
          end
          if(_zz_2[3100]) begin
            regVec_3100 <= _zz_regVec_0_1;
          end
          if(_zz_2[3101]) begin
            regVec_3101 <= _zz_regVec_0_1;
          end
          if(_zz_2[3102]) begin
            regVec_3102 <= _zz_regVec_0_1;
          end
          if(_zz_2[3103]) begin
            regVec_3103 <= _zz_regVec_0_1;
          end
          if(_zz_2[3104]) begin
            regVec_3104 <= _zz_regVec_0_1;
          end
          if(_zz_2[3105]) begin
            regVec_3105 <= _zz_regVec_0_1;
          end
          if(_zz_2[3106]) begin
            regVec_3106 <= _zz_regVec_0_1;
          end
          if(_zz_2[3107]) begin
            regVec_3107 <= _zz_regVec_0_1;
          end
          if(_zz_2[3108]) begin
            regVec_3108 <= _zz_regVec_0_1;
          end
          if(_zz_2[3109]) begin
            regVec_3109 <= _zz_regVec_0_1;
          end
          if(_zz_2[3110]) begin
            regVec_3110 <= _zz_regVec_0_1;
          end
          if(_zz_2[3111]) begin
            regVec_3111 <= _zz_regVec_0_1;
          end
          if(_zz_2[3112]) begin
            regVec_3112 <= _zz_regVec_0_1;
          end
          if(_zz_2[3113]) begin
            regVec_3113 <= _zz_regVec_0_1;
          end
          if(_zz_2[3114]) begin
            regVec_3114 <= _zz_regVec_0_1;
          end
          if(_zz_2[3115]) begin
            regVec_3115 <= _zz_regVec_0_1;
          end
          if(_zz_2[3116]) begin
            regVec_3116 <= _zz_regVec_0_1;
          end
          if(_zz_2[3117]) begin
            regVec_3117 <= _zz_regVec_0_1;
          end
          if(_zz_2[3118]) begin
            regVec_3118 <= _zz_regVec_0_1;
          end
          if(_zz_2[3119]) begin
            regVec_3119 <= _zz_regVec_0_1;
          end
          if(_zz_2[3120]) begin
            regVec_3120 <= _zz_regVec_0_1;
          end
          if(_zz_2[3121]) begin
            regVec_3121 <= _zz_regVec_0_1;
          end
          if(_zz_2[3122]) begin
            regVec_3122 <= _zz_regVec_0_1;
          end
          if(_zz_2[3123]) begin
            regVec_3123 <= _zz_regVec_0_1;
          end
          if(_zz_2[3124]) begin
            regVec_3124 <= _zz_regVec_0_1;
          end
          if(_zz_2[3125]) begin
            regVec_3125 <= _zz_regVec_0_1;
          end
          if(_zz_2[3126]) begin
            regVec_3126 <= _zz_regVec_0_1;
          end
          if(_zz_2[3127]) begin
            regVec_3127 <= _zz_regVec_0_1;
          end
          if(_zz_2[3128]) begin
            regVec_3128 <= _zz_regVec_0_1;
          end
          if(_zz_2[3129]) begin
            regVec_3129 <= _zz_regVec_0_1;
          end
          if(_zz_2[3130]) begin
            regVec_3130 <= _zz_regVec_0_1;
          end
          if(_zz_2[3131]) begin
            regVec_3131 <= _zz_regVec_0_1;
          end
          if(_zz_2[3132]) begin
            regVec_3132 <= _zz_regVec_0_1;
          end
          if(_zz_2[3133]) begin
            regVec_3133 <= _zz_regVec_0_1;
          end
          if(_zz_2[3134]) begin
            regVec_3134 <= _zz_regVec_0_1;
          end
          if(_zz_2[3135]) begin
            regVec_3135 <= _zz_regVec_0_1;
          end
          if(_zz_2[3136]) begin
            regVec_3136 <= _zz_regVec_0_1;
          end
          if(_zz_2[3137]) begin
            regVec_3137 <= _zz_regVec_0_1;
          end
          if(_zz_2[3138]) begin
            regVec_3138 <= _zz_regVec_0_1;
          end
          if(_zz_2[3139]) begin
            regVec_3139 <= _zz_regVec_0_1;
          end
          if(_zz_2[3140]) begin
            regVec_3140 <= _zz_regVec_0_1;
          end
          if(_zz_2[3141]) begin
            regVec_3141 <= _zz_regVec_0_1;
          end
          if(_zz_2[3142]) begin
            regVec_3142 <= _zz_regVec_0_1;
          end
          if(_zz_2[3143]) begin
            regVec_3143 <= _zz_regVec_0_1;
          end
          if(_zz_2[3144]) begin
            regVec_3144 <= _zz_regVec_0_1;
          end
          if(_zz_2[3145]) begin
            regVec_3145 <= _zz_regVec_0_1;
          end
          if(_zz_2[3146]) begin
            regVec_3146 <= _zz_regVec_0_1;
          end
          if(_zz_2[3147]) begin
            regVec_3147 <= _zz_regVec_0_1;
          end
          if(_zz_2[3148]) begin
            regVec_3148 <= _zz_regVec_0_1;
          end
          if(_zz_2[3149]) begin
            regVec_3149 <= _zz_regVec_0_1;
          end
          if(_zz_2[3150]) begin
            regVec_3150 <= _zz_regVec_0_1;
          end
          if(_zz_2[3151]) begin
            regVec_3151 <= _zz_regVec_0_1;
          end
          if(_zz_2[3152]) begin
            regVec_3152 <= _zz_regVec_0_1;
          end
          if(_zz_2[3153]) begin
            regVec_3153 <= _zz_regVec_0_1;
          end
          if(_zz_2[3154]) begin
            regVec_3154 <= _zz_regVec_0_1;
          end
          if(_zz_2[3155]) begin
            regVec_3155 <= _zz_regVec_0_1;
          end
          if(_zz_2[3156]) begin
            regVec_3156 <= _zz_regVec_0_1;
          end
          if(_zz_2[3157]) begin
            regVec_3157 <= _zz_regVec_0_1;
          end
          if(_zz_2[3158]) begin
            regVec_3158 <= _zz_regVec_0_1;
          end
          if(_zz_2[3159]) begin
            regVec_3159 <= _zz_regVec_0_1;
          end
          if(_zz_2[3160]) begin
            regVec_3160 <= _zz_regVec_0_1;
          end
          if(_zz_2[3161]) begin
            regVec_3161 <= _zz_regVec_0_1;
          end
          if(_zz_2[3162]) begin
            regVec_3162 <= _zz_regVec_0_1;
          end
          if(_zz_2[3163]) begin
            regVec_3163 <= _zz_regVec_0_1;
          end
          if(_zz_2[3164]) begin
            regVec_3164 <= _zz_regVec_0_1;
          end
          if(_zz_2[3165]) begin
            regVec_3165 <= _zz_regVec_0_1;
          end
          if(_zz_2[3166]) begin
            regVec_3166 <= _zz_regVec_0_1;
          end
          if(_zz_2[3167]) begin
            regVec_3167 <= _zz_regVec_0_1;
          end
          if(_zz_2[3168]) begin
            regVec_3168 <= _zz_regVec_0_1;
          end
          if(_zz_2[3169]) begin
            regVec_3169 <= _zz_regVec_0_1;
          end
          if(_zz_2[3170]) begin
            regVec_3170 <= _zz_regVec_0_1;
          end
          if(_zz_2[3171]) begin
            regVec_3171 <= _zz_regVec_0_1;
          end
          if(_zz_2[3172]) begin
            regVec_3172 <= _zz_regVec_0_1;
          end
          if(_zz_2[3173]) begin
            regVec_3173 <= _zz_regVec_0_1;
          end
          if(_zz_2[3174]) begin
            regVec_3174 <= _zz_regVec_0_1;
          end
          if(_zz_2[3175]) begin
            regVec_3175 <= _zz_regVec_0_1;
          end
          if(_zz_2[3176]) begin
            regVec_3176 <= _zz_regVec_0_1;
          end
          if(_zz_2[3177]) begin
            regVec_3177 <= _zz_regVec_0_1;
          end
          if(_zz_2[3178]) begin
            regVec_3178 <= _zz_regVec_0_1;
          end
          if(_zz_2[3179]) begin
            regVec_3179 <= _zz_regVec_0_1;
          end
          if(_zz_2[3180]) begin
            regVec_3180 <= _zz_regVec_0_1;
          end
          if(_zz_2[3181]) begin
            regVec_3181 <= _zz_regVec_0_1;
          end
          if(_zz_2[3182]) begin
            regVec_3182 <= _zz_regVec_0_1;
          end
          if(_zz_2[3183]) begin
            regVec_3183 <= _zz_regVec_0_1;
          end
          if(_zz_2[3184]) begin
            regVec_3184 <= _zz_regVec_0_1;
          end
          if(_zz_2[3185]) begin
            regVec_3185 <= _zz_regVec_0_1;
          end
          if(_zz_2[3186]) begin
            regVec_3186 <= _zz_regVec_0_1;
          end
          if(_zz_2[3187]) begin
            regVec_3187 <= _zz_regVec_0_1;
          end
          if(_zz_2[3188]) begin
            regVec_3188 <= _zz_regVec_0_1;
          end
          if(_zz_2[3189]) begin
            regVec_3189 <= _zz_regVec_0_1;
          end
          if(_zz_2[3190]) begin
            regVec_3190 <= _zz_regVec_0_1;
          end
          if(_zz_2[3191]) begin
            regVec_3191 <= _zz_regVec_0_1;
          end
          if(_zz_2[3192]) begin
            regVec_3192 <= _zz_regVec_0_1;
          end
          if(_zz_2[3193]) begin
            regVec_3193 <= _zz_regVec_0_1;
          end
          if(_zz_2[3194]) begin
            regVec_3194 <= _zz_regVec_0_1;
          end
          if(_zz_2[3195]) begin
            regVec_3195 <= _zz_regVec_0_1;
          end
          if(_zz_2[3196]) begin
            regVec_3196 <= _zz_regVec_0_1;
          end
          if(_zz_2[3197]) begin
            regVec_3197 <= _zz_regVec_0_1;
          end
          if(_zz_2[3198]) begin
            regVec_3198 <= _zz_regVec_0_1;
          end
          if(_zz_2[3199]) begin
            regVec_3199 <= _zz_regVec_0_1;
          end
          if(_zz_2[3200]) begin
            regVec_3200 <= _zz_regVec_0_1;
          end
          if(_zz_2[3201]) begin
            regVec_3201 <= _zz_regVec_0_1;
          end
          if(_zz_2[3202]) begin
            regVec_3202 <= _zz_regVec_0_1;
          end
          if(_zz_2[3203]) begin
            regVec_3203 <= _zz_regVec_0_1;
          end
          if(_zz_2[3204]) begin
            regVec_3204 <= _zz_regVec_0_1;
          end
          if(_zz_2[3205]) begin
            regVec_3205 <= _zz_regVec_0_1;
          end
          if(_zz_2[3206]) begin
            regVec_3206 <= _zz_regVec_0_1;
          end
          if(_zz_2[3207]) begin
            regVec_3207 <= _zz_regVec_0_1;
          end
          if(_zz_2[3208]) begin
            regVec_3208 <= _zz_regVec_0_1;
          end
          if(_zz_2[3209]) begin
            regVec_3209 <= _zz_regVec_0_1;
          end
          if(_zz_2[3210]) begin
            regVec_3210 <= _zz_regVec_0_1;
          end
          if(_zz_2[3211]) begin
            regVec_3211 <= _zz_regVec_0_1;
          end
          if(_zz_2[3212]) begin
            regVec_3212 <= _zz_regVec_0_1;
          end
          if(_zz_2[3213]) begin
            regVec_3213 <= _zz_regVec_0_1;
          end
          if(_zz_2[3214]) begin
            regVec_3214 <= _zz_regVec_0_1;
          end
          if(_zz_2[3215]) begin
            regVec_3215 <= _zz_regVec_0_1;
          end
          if(_zz_2[3216]) begin
            regVec_3216 <= _zz_regVec_0_1;
          end
          if(_zz_2[3217]) begin
            regVec_3217 <= _zz_regVec_0_1;
          end
          if(_zz_2[3218]) begin
            regVec_3218 <= _zz_regVec_0_1;
          end
          if(_zz_2[3219]) begin
            regVec_3219 <= _zz_regVec_0_1;
          end
          if(_zz_2[3220]) begin
            regVec_3220 <= _zz_regVec_0_1;
          end
          if(_zz_2[3221]) begin
            regVec_3221 <= _zz_regVec_0_1;
          end
          if(_zz_2[3222]) begin
            regVec_3222 <= _zz_regVec_0_1;
          end
          if(_zz_2[3223]) begin
            regVec_3223 <= _zz_regVec_0_1;
          end
          if(_zz_2[3224]) begin
            regVec_3224 <= _zz_regVec_0_1;
          end
          if(_zz_2[3225]) begin
            regVec_3225 <= _zz_regVec_0_1;
          end
          if(_zz_2[3226]) begin
            regVec_3226 <= _zz_regVec_0_1;
          end
          if(_zz_2[3227]) begin
            regVec_3227 <= _zz_regVec_0_1;
          end
          if(_zz_2[3228]) begin
            regVec_3228 <= _zz_regVec_0_1;
          end
          if(_zz_2[3229]) begin
            regVec_3229 <= _zz_regVec_0_1;
          end
          if(_zz_2[3230]) begin
            regVec_3230 <= _zz_regVec_0_1;
          end
          if(_zz_2[3231]) begin
            regVec_3231 <= _zz_regVec_0_1;
          end
          if(_zz_2[3232]) begin
            regVec_3232 <= _zz_regVec_0_1;
          end
          if(_zz_2[3233]) begin
            regVec_3233 <= _zz_regVec_0_1;
          end
          if(_zz_2[3234]) begin
            regVec_3234 <= _zz_regVec_0_1;
          end
          if(_zz_2[3235]) begin
            regVec_3235 <= _zz_regVec_0_1;
          end
          if(_zz_2[3236]) begin
            regVec_3236 <= _zz_regVec_0_1;
          end
          if(_zz_2[3237]) begin
            regVec_3237 <= _zz_regVec_0_1;
          end
          if(_zz_2[3238]) begin
            regVec_3238 <= _zz_regVec_0_1;
          end
          if(_zz_2[3239]) begin
            regVec_3239 <= _zz_regVec_0_1;
          end
          if(_zz_2[3240]) begin
            regVec_3240 <= _zz_regVec_0_1;
          end
          if(_zz_2[3241]) begin
            regVec_3241 <= _zz_regVec_0_1;
          end
          if(_zz_2[3242]) begin
            regVec_3242 <= _zz_regVec_0_1;
          end
          if(_zz_2[3243]) begin
            regVec_3243 <= _zz_regVec_0_1;
          end
          if(_zz_2[3244]) begin
            regVec_3244 <= _zz_regVec_0_1;
          end
          if(_zz_2[3245]) begin
            regVec_3245 <= _zz_regVec_0_1;
          end
          if(_zz_2[3246]) begin
            regVec_3246 <= _zz_regVec_0_1;
          end
          if(_zz_2[3247]) begin
            regVec_3247 <= _zz_regVec_0_1;
          end
          if(_zz_2[3248]) begin
            regVec_3248 <= _zz_regVec_0_1;
          end
          if(_zz_2[3249]) begin
            regVec_3249 <= _zz_regVec_0_1;
          end
          if(_zz_2[3250]) begin
            regVec_3250 <= _zz_regVec_0_1;
          end
          if(_zz_2[3251]) begin
            regVec_3251 <= _zz_regVec_0_1;
          end
          if(_zz_2[3252]) begin
            regVec_3252 <= _zz_regVec_0_1;
          end
          if(_zz_2[3253]) begin
            regVec_3253 <= _zz_regVec_0_1;
          end
          if(_zz_2[3254]) begin
            regVec_3254 <= _zz_regVec_0_1;
          end
          if(_zz_2[3255]) begin
            regVec_3255 <= _zz_regVec_0_1;
          end
          if(_zz_2[3256]) begin
            regVec_3256 <= _zz_regVec_0_1;
          end
          if(_zz_2[3257]) begin
            regVec_3257 <= _zz_regVec_0_1;
          end
          if(_zz_2[3258]) begin
            regVec_3258 <= _zz_regVec_0_1;
          end
          if(_zz_2[3259]) begin
            regVec_3259 <= _zz_regVec_0_1;
          end
          if(_zz_2[3260]) begin
            regVec_3260 <= _zz_regVec_0_1;
          end
          if(_zz_2[3261]) begin
            regVec_3261 <= _zz_regVec_0_1;
          end
          if(_zz_2[3262]) begin
            regVec_3262 <= _zz_regVec_0_1;
          end
          if(_zz_2[3263]) begin
            regVec_3263 <= _zz_regVec_0_1;
          end
          if(_zz_2[3264]) begin
            regVec_3264 <= _zz_regVec_0_1;
          end
          if(_zz_2[3265]) begin
            regVec_3265 <= _zz_regVec_0_1;
          end
          if(_zz_2[3266]) begin
            regVec_3266 <= _zz_regVec_0_1;
          end
          if(_zz_2[3267]) begin
            regVec_3267 <= _zz_regVec_0_1;
          end
          if(_zz_2[3268]) begin
            regVec_3268 <= _zz_regVec_0_1;
          end
          if(_zz_2[3269]) begin
            regVec_3269 <= _zz_regVec_0_1;
          end
          if(_zz_2[3270]) begin
            regVec_3270 <= _zz_regVec_0_1;
          end
          if(_zz_2[3271]) begin
            regVec_3271 <= _zz_regVec_0_1;
          end
          if(_zz_2[3272]) begin
            regVec_3272 <= _zz_regVec_0_1;
          end
          if(_zz_2[3273]) begin
            regVec_3273 <= _zz_regVec_0_1;
          end
          if(_zz_2[3274]) begin
            regVec_3274 <= _zz_regVec_0_1;
          end
          if(_zz_2[3275]) begin
            regVec_3275 <= _zz_regVec_0_1;
          end
          if(_zz_2[3276]) begin
            regVec_3276 <= _zz_regVec_0_1;
          end
          if(_zz_2[3277]) begin
            regVec_3277 <= _zz_regVec_0_1;
          end
          if(_zz_2[3278]) begin
            regVec_3278 <= _zz_regVec_0_1;
          end
          if(_zz_2[3279]) begin
            regVec_3279 <= _zz_regVec_0_1;
          end
          if(_zz_2[3280]) begin
            regVec_3280 <= _zz_regVec_0_1;
          end
          if(_zz_2[3281]) begin
            regVec_3281 <= _zz_regVec_0_1;
          end
          if(_zz_2[3282]) begin
            regVec_3282 <= _zz_regVec_0_1;
          end
          if(_zz_2[3283]) begin
            regVec_3283 <= _zz_regVec_0_1;
          end
          if(_zz_2[3284]) begin
            regVec_3284 <= _zz_regVec_0_1;
          end
          if(_zz_2[3285]) begin
            regVec_3285 <= _zz_regVec_0_1;
          end
          if(_zz_2[3286]) begin
            regVec_3286 <= _zz_regVec_0_1;
          end
          if(_zz_2[3287]) begin
            regVec_3287 <= _zz_regVec_0_1;
          end
          if(_zz_2[3288]) begin
            regVec_3288 <= _zz_regVec_0_1;
          end
          if(_zz_2[3289]) begin
            regVec_3289 <= _zz_regVec_0_1;
          end
          if(_zz_2[3290]) begin
            regVec_3290 <= _zz_regVec_0_1;
          end
          if(_zz_2[3291]) begin
            regVec_3291 <= _zz_regVec_0_1;
          end
          if(_zz_2[3292]) begin
            regVec_3292 <= _zz_regVec_0_1;
          end
          if(_zz_2[3293]) begin
            regVec_3293 <= _zz_regVec_0_1;
          end
          if(_zz_2[3294]) begin
            regVec_3294 <= _zz_regVec_0_1;
          end
          if(_zz_2[3295]) begin
            regVec_3295 <= _zz_regVec_0_1;
          end
          if(_zz_2[3296]) begin
            regVec_3296 <= _zz_regVec_0_1;
          end
          if(_zz_2[3297]) begin
            regVec_3297 <= _zz_regVec_0_1;
          end
          if(_zz_2[3298]) begin
            regVec_3298 <= _zz_regVec_0_1;
          end
          if(_zz_2[3299]) begin
            regVec_3299 <= _zz_regVec_0_1;
          end
          if(_zz_2[3300]) begin
            regVec_3300 <= _zz_regVec_0_1;
          end
          if(_zz_2[3301]) begin
            regVec_3301 <= _zz_regVec_0_1;
          end
          if(_zz_2[3302]) begin
            regVec_3302 <= _zz_regVec_0_1;
          end
          if(_zz_2[3303]) begin
            regVec_3303 <= _zz_regVec_0_1;
          end
          if(_zz_2[3304]) begin
            regVec_3304 <= _zz_regVec_0_1;
          end
          if(_zz_2[3305]) begin
            regVec_3305 <= _zz_regVec_0_1;
          end
          if(_zz_2[3306]) begin
            regVec_3306 <= _zz_regVec_0_1;
          end
          if(_zz_2[3307]) begin
            regVec_3307 <= _zz_regVec_0_1;
          end
          if(_zz_2[3308]) begin
            regVec_3308 <= _zz_regVec_0_1;
          end
          if(_zz_2[3309]) begin
            regVec_3309 <= _zz_regVec_0_1;
          end
          if(_zz_2[3310]) begin
            regVec_3310 <= _zz_regVec_0_1;
          end
          if(_zz_2[3311]) begin
            regVec_3311 <= _zz_regVec_0_1;
          end
          if(_zz_2[3312]) begin
            regVec_3312 <= _zz_regVec_0_1;
          end
          if(_zz_2[3313]) begin
            regVec_3313 <= _zz_regVec_0_1;
          end
          if(_zz_2[3314]) begin
            regVec_3314 <= _zz_regVec_0_1;
          end
          if(_zz_2[3315]) begin
            regVec_3315 <= _zz_regVec_0_1;
          end
          if(_zz_2[3316]) begin
            regVec_3316 <= _zz_regVec_0_1;
          end
          if(_zz_2[3317]) begin
            regVec_3317 <= _zz_regVec_0_1;
          end
          if(_zz_2[3318]) begin
            regVec_3318 <= _zz_regVec_0_1;
          end
          if(_zz_2[3319]) begin
            regVec_3319 <= _zz_regVec_0_1;
          end
          if(_zz_2[3320]) begin
            regVec_3320 <= _zz_regVec_0_1;
          end
          if(_zz_2[3321]) begin
            regVec_3321 <= _zz_regVec_0_1;
          end
          if(_zz_2[3322]) begin
            regVec_3322 <= _zz_regVec_0_1;
          end
          if(_zz_2[3323]) begin
            regVec_3323 <= _zz_regVec_0_1;
          end
          if(_zz_2[3324]) begin
            regVec_3324 <= _zz_regVec_0_1;
          end
          if(_zz_2[3325]) begin
            regVec_3325 <= _zz_regVec_0_1;
          end
          if(_zz_2[3326]) begin
            regVec_3326 <= _zz_regVec_0_1;
          end
          if(_zz_2[3327]) begin
            regVec_3327 <= _zz_regVec_0_1;
          end
          if(_zz_2[3328]) begin
            regVec_3328 <= _zz_regVec_0_1;
          end
          if(_zz_2[3329]) begin
            regVec_3329 <= _zz_regVec_0_1;
          end
          if(_zz_2[3330]) begin
            regVec_3330 <= _zz_regVec_0_1;
          end
          if(_zz_2[3331]) begin
            regVec_3331 <= _zz_regVec_0_1;
          end
          if(_zz_2[3332]) begin
            regVec_3332 <= _zz_regVec_0_1;
          end
          if(_zz_2[3333]) begin
            regVec_3333 <= _zz_regVec_0_1;
          end
          if(_zz_2[3334]) begin
            regVec_3334 <= _zz_regVec_0_1;
          end
          if(_zz_2[3335]) begin
            regVec_3335 <= _zz_regVec_0_1;
          end
          if(_zz_2[3336]) begin
            regVec_3336 <= _zz_regVec_0_1;
          end
          if(_zz_2[3337]) begin
            regVec_3337 <= _zz_regVec_0_1;
          end
          if(_zz_2[3338]) begin
            regVec_3338 <= _zz_regVec_0_1;
          end
          if(_zz_2[3339]) begin
            regVec_3339 <= _zz_regVec_0_1;
          end
          if(_zz_2[3340]) begin
            regVec_3340 <= _zz_regVec_0_1;
          end
          if(_zz_2[3341]) begin
            regVec_3341 <= _zz_regVec_0_1;
          end
          if(_zz_2[3342]) begin
            regVec_3342 <= _zz_regVec_0_1;
          end
          if(_zz_2[3343]) begin
            regVec_3343 <= _zz_regVec_0_1;
          end
          if(_zz_2[3344]) begin
            regVec_3344 <= _zz_regVec_0_1;
          end
          if(_zz_2[3345]) begin
            regVec_3345 <= _zz_regVec_0_1;
          end
          if(_zz_2[3346]) begin
            regVec_3346 <= _zz_regVec_0_1;
          end
          if(_zz_2[3347]) begin
            regVec_3347 <= _zz_regVec_0_1;
          end
          if(_zz_2[3348]) begin
            regVec_3348 <= _zz_regVec_0_1;
          end
          if(_zz_2[3349]) begin
            regVec_3349 <= _zz_regVec_0_1;
          end
          if(_zz_2[3350]) begin
            regVec_3350 <= _zz_regVec_0_1;
          end
          if(_zz_2[3351]) begin
            regVec_3351 <= _zz_regVec_0_1;
          end
          if(_zz_2[3352]) begin
            regVec_3352 <= _zz_regVec_0_1;
          end
          if(_zz_2[3353]) begin
            regVec_3353 <= _zz_regVec_0_1;
          end
          if(_zz_2[3354]) begin
            regVec_3354 <= _zz_regVec_0_1;
          end
          if(_zz_2[3355]) begin
            regVec_3355 <= _zz_regVec_0_1;
          end
          if(_zz_2[3356]) begin
            regVec_3356 <= _zz_regVec_0_1;
          end
          if(_zz_2[3357]) begin
            regVec_3357 <= _zz_regVec_0_1;
          end
          if(_zz_2[3358]) begin
            regVec_3358 <= _zz_regVec_0_1;
          end
          if(_zz_2[3359]) begin
            regVec_3359 <= _zz_regVec_0_1;
          end
          if(_zz_2[3360]) begin
            regVec_3360 <= _zz_regVec_0_1;
          end
          if(_zz_2[3361]) begin
            regVec_3361 <= _zz_regVec_0_1;
          end
          if(_zz_2[3362]) begin
            regVec_3362 <= _zz_regVec_0_1;
          end
          if(_zz_2[3363]) begin
            regVec_3363 <= _zz_regVec_0_1;
          end
          if(_zz_2[3364]) begin
            regVec_3364 <= _zz_regVec_0_1;
          end
          if(_zz_2[3365]) begin
            regVec_3365 <= _zz_regVec_0_1;
          end
          if(_zz_2[3366]) begin
            regVec_3366 <= _zz_regVec_0_1;
          end
          if(_zz_2[3367]) begin
            regVec_3367 <= _zz_regVec_0_1;
          end
          if(_zz_2[3368]) begin
            regVec_3368 <= _zz_regVec_0_1;
          end
          if(_zz_2[3369]) begin
            regVec_3369 <= _zz_regVec_0_1;
          end
          if(_zz_2[3370]) begin
            regVec_3370 <= _zz_regVec_0_1;
          end
          if(_zz_2[3371]) begin
            regVec_3371 <= _zz_regVec_0_1;
          end
          if(_zz_2[3372]) begin
            regVec_3372 <= _zz_regVec_0_1;
          end
          if(_zz_2[3373]) begin
            regVec_3373 <= _zz_regVec_0_1;
          end
          if(_zz_2[3374]) begin
            regVec_3374 <= _zz_regVec_0_1;
          end
          if(_zz_2[3375]) begin
            regVec_3375 <= _zz_regVec_0_1;
          end
          if(_zz_2[3376]) begin
            regVec_3376 <= _zz_regVec_0_1;
          end
          if(_zz_2[3377]) begin
            regVec_3377 <= _zz_regVec_0_1;
          end
          if(_zz_2[3378]) begin
            regVec_3378 <= _zz_regVec_0_1;
          end
          if(_zz_2[3379]) begin
            regVec_3379 <= _zz_regVec_0_1;
          end
          if(_zz_2[3380]) begin
            regVec_3380 <= _zz_regVec_0_1;
          end
          if(_zz_2[3381]) begin
            regVec_3381 <= _zz_regVec_0_1;
          end
          if(_zz_2[3382]) begin
            regVec_3382 <= _zz_regVec_0_1;
          end
          if(_zz_2[3383]) begin
            regVec_3383 <= _zz_regVec_0_1;
          end
          if(_zz_2[3384]) begin
            regVec_3384 <= _zz_regVec_0_1;
          end
          if(_zz_2[3385]) begin
            regVec_3385 <= _zz_regVec_0_1;
          end
          if(_zz_2[3386]) begin
            regVec_3386 <= _zz_regVec_0_1;
          end
          if(_zz_2[3387]) begin
            regVec_3387 <= _zz_regVec_0_1;
          end
          if(_zz_2[3388]) begin
            regVec_3388 <= _zz_regVec_0_1;
          end
          if(_zz_2[3389]) begin
            regVec_3389 <= _zz_regVec_0_1;
          end
          if(_zz_2[3390]) begin
            regVec_3390 <= _zz_regVec_0_1;
          end
          if(_zz_2[3391]) begin
            regVec_3391 <= _zz_regVec_0_1;
          end
          if(_zz_2[3392]) begin
            regVec_3392 <= _zz_regVec_0_1;
          end
          if(_zz_2[3393]) begin
            regVec_3393 <= _zz_regVec_0_1;
          end
          if(_zz_2[3394]) begin
            regVec_3394 <= _zz_regVec_0_1;
          end
          if(_zz_2[3395]) begin
            regVec_3395 <= _zz_regVec_0_1;
          end
          if(_zz_2[3396]) begin
            regVec_3396 <= _zz_regVec_0_1;
          end
          if(_zz_2[3397]) begin
            regVec_3397 <= _zz_regVec_0_1;
          end
          if(_zz_2[3398]) begin
            regVec_3398 <= _zz_regVec_0_1;
          end
          if(_zz_2[3399]) begin
            regVec_3399 <= _zz_regVec_0_1;
          end
          if(_zz_2[3400]) begin
            regVec_3400 <= _zz_regVec_0_1;
          end
          if(_zz_2[3401]) begin
            regVec_3401 <= _zz_regVec_0_1;
          end
          if(_zz_2[3402]) begin
            regVec_3402 <= _zz_regVec_0_1;
          end
          if(_zz_2[3403]) begin
            regVec_3403 <= _zz_regVec_0_1;
          end
          if(_zz_2[3404]) begin
            regVec_3404 <= _zz_regVec_0_1;
          end
          if(_zz_2[3405]) begin
            regVec_3405 <= _zz_regVec_0_1;
          end
          if(_zz_2[3406]) begin
            regVec_3406 <= _zz_regVec_0_1;
          end
          if(_zz_2[3407]) begin
            regVec_3407 <= _zz_regVec_0_1;
          end
          if(_zz_2[3408]) begin
            regVec_3408 <= _zz_regVec_0_1;
          end
          if(_zz_2[3409]) begin
            regVec_3409 <= _zz_regVec_0_1;
          end
          if(_zz_2[3410]) begin
            regVec_3410 <= _zz_regVec_0_1;
          end
          if(_zz_2[3411]) begin
            regVec_3411 <= _zz_regVec_0_1;
          end
          if(_zz_2[3412]) begin
            regVec_3412 <= _zz_regVec_0_1;
          end
          if(_zz_2[3413]) begin
            regVec_3413 <= _zz_regVec_0_1;
          end
          if(_zz_2[3414]) begin
            regVec_3414 <= _zz_regVec_0_1;
          end
          if(_zz_2[3415]) begin
            regVec_3415 <= _zz_regVec_0_1;
          end
          if(_zz_2[3416]) begin
            regVec_3416 <= _zz_regVec_0_1;
          end
          if(_zz_2[3417]) begin
            regVec_3417 <= _zz_regVec_0_1;
          end
          if(_zz_2[3418]) begin
            regVec_3418 <= _zz_regVec_0_1;
          end
          if(_zz_2[3419]) begin
            regVec_3419 <= _zz_regVec_0_1;
          end
          if(_zz_2[3420]) begin
            regVec_3420 <= _zz_regVec_0_1;
          end
          if(_zz_2[3421]) begin
            regVec_3421 <= _zz_regVec_0_1;
          end
          if(_zz_2[3422]) begin
            regVec_3422 <= _zz_regVec_0_1;
          end
          if(_zz_2[3423]) begin
            regVec_3423 <= _zz_regVec_0_1;
          end
          if(_zz_2[3424]) begin
            regVec_3424 <= _zz_regVec_0_1;
          end
          if(_zz_2[3425]) begin
            regVec_3425 <= _zz_regVec_0_1;
          end
          if(_zz_2[3426]) begin
            regVec_3426 <= _zz_regVec_0_1;
          end
          if(_zz_2[3427]) begin
            regVec_3427 <= _zz_regVec_0_1;
          end
          if(_zz_2[3428]) begin
            regVec_3428 <= _zz_regVec_0_1;
          end
          if(_zz_2[3429]) begin
            regVec_3429 <= _zz_regVec_0_1;
          end
          if(_zz_2[3430]) begin
            regVec_3430 <= _zz_regVec_0_1;
          end
          if(_zz_2[3431]) begin
            regVec_3431 <= _zz_regVec_0_1;
          end
          if(_zz_2[3432]) begin
            regVec_3432 <= _zz_regVec_0_1;
          end
          if(_zz_2[3433]) begin
            regVec_3433 <= _zz_regVec_0_1;
          end
          if(_zz_2[3434]) begin
            regVec_3434 <= _zz_regVec_0_1;
          end
          if(_zz_2[3435]) begin
            regVec_3435 <= _zz_regVec_0_1;
          end
          if(_zz_2[3436]) begin
            regVec_3436 <= _zz_regVec_0_1;
          end
          if(_zz_2[3437]) begin
            regVec_3437 <= _zz_regVec_0_1;
          end
          if(_zz_2[3438]) begin
            regVec_3438 <= _zz_regVec_0_1;
          end
          if(_zz_2[3439]) begin
            regVec_3439 <= _zz_regVec_0_1;
          end
          if(_zz_2[3440]) begin
            regVec_3440 <= _zz_regVec_0_1;
          end
          if(_zz_2[3441]) begin
            regVec_3441 <= _zz_regVec_0_1;
          end
          if(_zz_2[3442]) begin
            regVec_3442 <= _zz_regVec_0_1;
          end
          if(_zz_2[3443]) begin
            regVec_3443 <= _zz_regVec_0_1;
          end
          if(_zz_2[3444]) begin
            regVec_3444 <= _zz_regVec_0_1;
          end
          if(_zz_2[3445]) begin
            regVec_3445 <= _zz_regVec_0_1;
          end
          if(_zz_2[3446]) begin
            regVec_3446 <= _zz_regVec_0_1;
          end
          if(_zz_2[3447]) begin
            regVec_3447 <= _zz_regVec_0_1;
          end
          if(_zz_2[3448]) begin
            regVec_3448 <= _zz_regVec_0_1;
          end
          if(_zz_2[3449]) begin
            regVec_3449 <= _zz_regVec_0_1;
          end
          if(_zz_2[3450]) begin
            regVec_3450 <= _zz_regVec_0_1;
          end
          if(_zz_2[3451]) begin
            regVec_3451 <= _zz_regVec_0_1;
          end
          if(_zz_2[3452]) begin
            regVec_3452 <= _zz_regVec_0_1;
          end
          if(_zz_2[3453]) begin
            regVec_3453 <= _zz_regVec_0_1;
          end
          if(_zz_2[3454]) begin
            regVec_3454 <= _zz_regVec_0_1;
          end
          if(_zz_2[3455]) begin
            regVec_3455 <= _zz_regVec_0_1;
          end
          if(_zz_2[3456]) begin
            regVec_3456 <= _zz_regVec_0_1;
          end
          if(_zz_2[3457]) begin
            regVec_3457 <= _zz_regVec_0_1;
          end
          if(_zz_2[3458]) begin
            regVec_3458 <= _zz_regVec_0_1;
          end
          if(_zz_2[3459]) begin
            regVec_3459 <= _zz_regVec_0_1;
          end
          if(_zz_2[3460]) begin
            regVec_3460 <= _zz_regVec_0_1;
          end
          if(_zz_2[3461]) begin
            regVec_3461 <= _zz_regVec_0_1;
          end
          if(_zz_2[3462]) begin
            regVec_3462 <= _zz_regVec_0_1;
          end
          if(_zz_2[3463]) begin
            regVec_3463 <= _zz_regVec_0_1;
          end
          if(_zz_2[3464]) begin
            regVec_3464 <= _zz_regVec_0_1;
          end
          if(_zz_2[3465]) begin
            regVec_3465 <= _zz_regVec_0_1;
          end
          if(_zz_2[3466]) begin
            regVec_3466 <= _zz_regVec_0_1;
          end
          if(_zz_2[3467]) begin
            regVec_3467 <= _zz_regVec_0_1;
          end
          if(_zz_2[3468]) begin
            regVec_3468 <= _zz_regVec_0_1;
          end
          if(_zz_2[3469]) begin
            regVec_3469 <= _zz_regVec_0_1;
          end
          if(_zz_2[3470]) begin
            regVec_3470 <= _zz_regVec_0_1;
          end
          if(_zz_2[3471]) begin
            regVec_3471 <= _zz_regVec_0_1;
          end
          if(_zz_2[3472]) begin
            regVec_3472 <= _zz_regVec_0_1;
          end
          if(_zz_2[3473]) begin
            regVec_3473 <= _zz_regVec_0_1;
          end
          if(_zz_2[3474]) begin
            regVec_3474 <= _zz_regVec_0_1;
          end
          if(_zz_2[3475]) begin
            regVec_3475 <= _zz_regVec_0_1;
          end
          if(_zz_2[3476]) begin
            regVec_3476 <= _zz_regVec_0_1;
          end
          if(_zz_2[3477]) begin
            regVec_3477 <= _zz_regVec_0_1;
          end
          if(_zz_2[3478]) begin
            regVec_3478 <= _zz_regVec_0_1;
          end
          if(_zz_2[3479]) begin
            regVec_3479 <= _zz_regVec_0_1;
          end
          if(_zz_2[3480]) begin
            regVec_3480 <= _zz_regVec_0_1;
          end
          if(_zz_2[3481]) begin
            regVec_3481 <= _zz_regVec_0_1;
          end
          if(_zz_2[3482]) begin
            regVec_3482 <= _zz_regVec_0_1;
          end
          if(_zz_2[3483]) begin
            regVec_3483 <= _zz_regVec_0_1;
          end
          if(_zz_2[3484]) begin
            regVec_3484 <= _zz_regVec_0_1;
          end
          if(_zz_2[3485]) begin
            regVec_3485 <= _zz_regVec_0_1;
          end
          if(_zz_2[3486]) begin
            regVec_3486 <= _zz_regVec_0_1;
          end
          if(_zz_2[3487]) begin
            regVec_3487 <= _zz_regVec_0_1;
          end
          if(_zz_2[3488]) begin
            regVec_3488 <= _zz_regVec_0_1;
          end
          if(_zz_2[3489]) begin
            regVec_3489 <= _zz_regVec_0_1;
          end
          if(_zz_2[3490]) begin
            regVec_3490 <= _zz_regVec_0_1;
          end
          if(_zz_2[3491]) begin
            regVec_3491 <= _zz_regVec_0_1;
          end
          if(_zz_2[3492]) begin
            regVec_3492 <= _zz_regVec_0_1;
          end
          if(_zz_2[3493]) begin
            regVec_3493 <= _zz_regVec_0_1;
          end
          if(_zz_2[3494]) begin
            regVec_3494 <= _zz_regVec_0_1;
          end
          if(_zz_2[3495]) begin
            regVec_3495 <= _zz_regVec_0_1;
          end
          if(_zz_2[3496]) begin
            regVec_3496 <= _zz_regVec_0_1;
          end
          if(_zz_2[3497]) begin
            regVec_3497 <= _zz_regVec_0_1;
          end
          if(_zz_2[3498]) begin
            regVec_3498 <= _zz_regVec_0_1;
          end
          if(_zz_2[3499]) begin
            regVec_3499 <= _zz_regVec_0_1;
          end
          if(_zz_2[3500]) begin
            regVec_3500 <= _zz_regVec_0_1;
          end
          if(_zz_2[3501]) begin
            regVec_3501 <= _zz_regVec_0_1;
          end
          if(_zz_2[3502]) begin
            regVec_3502 <= _zz_regVec_0_1;
          end
          if(_zz_2[3503]) begin
            regVec_3503 <= _zz_regVec_0_1;
          end
          if(_zz_2[3504]) begin
            regVec_3504 <= _zz_regVec_0_1;
          end
          if(_zz_2[3505]) begin
            regVec_3505 <= _zz_regVec_0_1;
          end
          if(_zz_2[3506]) begin
            regVec_3506 <= _zz_regVec_0_1;
          end
          if(_zz_2[3507]) begin
            regVec_3507 <= _zz_regVec_0_1;
          end
          if(_zz_2[3508]) begin
            regVec_3508 <= _zz_regVec_0_1;
          end
          if(_zz_2[3509]) begin
            regVec_3509 <= _zz_regVec_0_1;
          end
          if(_zz_2[3510]) begin
            regVec_3510 <= _zz_regVec_0_1;
          end
          if(_zz_2[3511]) begin
            regVec_3511 <= _zz_regVec_0_1;
          end
          if(_zz_2[3512]) begin
            regVec_3512 <= _zz_regVec_0_1;
          end
          if(_zz_2[3513]) begin
            regVec_3513 <= _zz_regVec_0_1;
          end
          if(_zz_2[3514]) begin
            regVec_3514 <= _zz_regVec_0_1;
          end
          if(_zz_2[3515]) begin
            regVec_3515 <= _zz_regVec_0_1;
          end
          if(_zz_2[3516]) begin
            regVec_3516 <= _zz_regVec_0_1;
          end
          if(_zz_2[3517]) begin
            regVec_3517 <= _zz_regVec_0_1;
          end
          if(_zz_2[3518]) begin
            regVec_3518 <= _zz_regVec_0_1;
          end
          if(_zz_2[3519]) begin
            regVec_3519 <= _zz_regVec_0_1;
          end
          if(_zz_2[3520]) begin
            regVec_3520 <= _zz_regVec_0_1;
          end
          if(_zz_2[3521]) begin
            regVec_3521 <= _zz_regVec_0_1;
          end
          if(_zz_2[3522]) begin
            regVec_3522 <= _zz_regVec_0_1;
          end
          if(_zz_2[3523]) begin
            regVec_3523 <= _zz_regVec_0_1;
          end
          if(_zz_2[3524]) begin
            regVec_3524 <= _zz_regVec_0_1;
          end
          if(_zz_2[3525]) begin
            regVec_3525 <= _zz_regVec_0_1;
          end
          if(_zz_2[3526]) begin
            regVec_3526 <= _zz_regVec_0_1;
          end
          if(_zz_2[3527]) begin
            regVec_3527 <= _zz_regVec_0_1;
          end
          if(_zz_2[3528]) begin
            regVec_3528 <= _zz_regVec_0_1;
          end
          if(_zz_2[3529]) begin
            regVec_3529 <= _zz_regVec_0_1;
          end
          if(_zz_2[3530]) begin
            regVec_3530 <= _zz_regVec_0_1;
          end
          if(_zz_2[3531]) begin
            regVec_3531 <= _zz_regVec_0_1;
          end
          if(_zz_2[3532]) begin
            regVec_3532 <= _zz_regVec_0_1;
          end
          if(_zz_2[3533]) begin
            regVec_3533 <= _zz_regVec_0_1;
          end
          if(_zz_2[3534]) begin
            regVec_3534 <= _zz_regVec_0_1;
          end
          if(_zz_2[3535]) begin
            regVec_3535 <= _zz_regVec_0_1;
          end
          if(_zz_2[3536]) begin
            regVec_3536 <= _zz_regVec_0_1;
          end
          if(_zz_2[3537]) begin
            regVec_3537 <= _zz_regVec_0_1;
          end
          if(_zz_2[3538]) begin
            regVec_3538 <= _zz_regVec_0_1;
          end
          if(_zz_2[3539]) begin
            regVec_3539 <= _zz_regVec_0_1;
          end
          if(_zz_2[3540]) begin
            regVec_3540 <= _zz_regVec_0_1;
          end
          if(_zz_2[3541]) begin
            regVec_3541 <= _zz_regVec_0_1;
          end
          if(_zz_2[3542]) begin
            regVec_3542 <= _zz_regVec_0_1;
          end
          if(_zz_2[3543]) begin
            regVec_3543 <= _zz_regVec_0_1;
          end
          if(_zz_2[3544]) begin
            regVec_3544 <= _zz_regVec_0_1;
          end
          if(_zz_2[3545]) begin
            regVec_3545 <= _zz_regVec_0_1;
          end
          if(_zz_2[3546]) begin
            regVec_3546 <= _zz_regVec_0_1;
          end
          if(_zz_2[3547]) begin
            regVec_3547 <= _zz_regVec_0_1;
          end
          if(_zz_2[3548]) begin
            regVec_3548 <= _zz_regVec_0_1;
          end
          if(_zz_2[3549]) begin
            regVec_3549 <= _zz_regVec_0_1;
          end
          if(_zz_2[3550]) begin
            regVec_3550 <= _zz_regVec_0_1;
          end
          if(_zz_2[3551]) begin
            regVec_3551 <= _zz_regVec_0_1;
          end
          if(_zz_2[3552]) begin
            regVec_3552 <= _zz_regVec_0_1;
          end
          if(_zz_2[3553]) begin
            regVec_3553 <= _zz_regVec_0_1;
          end
          if(_zz_2[3554]) begin
            regVec_3554 <= _zz_regVec_0_1;
          end
          if(_zz_2[3555]) begin
            regVec_3555 <= _zz_regVec_0_1;
          end
          if(_zz_2[3556]) begin
            regVec_3556 <= _zz_regVec_0_1;
          end
          if(_zz_2[3557]) begin
            regVec_3557 <= _zz_regVec_0_1;
          end
          if(_zz_2[3558]) begin
            regVec_3558 <= _zz_regVec_0_1;
          end
          if(_zz_2[3559]) begin
            regVec_3559 <= _zz_regVec_0_1;
          end
          if(_zz_2[3560]) begin
            regVec_3560 <= _zz_regVec_0_1;
          end
          if(_zz_2[3561]) begin
            regVec_3561 <= _zz_regVec_0_1;
          end
          if(_zz_2[3562]) begin
            regVec_3562 <= _zz_regVec_0_1;
          end
          if(_zz_2[3563]) begin
            regVec_3563 <= _zz_regVec_0_1;
          end
          if(_zz_2[3564]) begin
            regVec_3564 <= _zz_regVec_0_1;
          end
          if(_zz_2[3565]) begin
            regVec_3565 <= _zz_regVec_0_1;
          end
          if(_zz_2[3566]) begin
            regVec_3566 <= _zz_regVec_0_1;
          end
          if(_zz_2[3567]) begin
            regVec_3567 <= _zz_regVec_0_1;
          end
          if(_zz_2[3568]) begin
            regVec_3568 <= _zz_regVec_0_1;
          end
          if(_zz_2[3569]) begin
            regVec_3569 <= _zz_regVec_0_1;
          end
          if(_zz_2[3570]) begin
            regVec_3570 <= _zz_regVec_0_1;
          end
          if(_zz_2[3571]) begin
            regVec_3571 <= _zz_regVec_0_1;
          end
          if(_zz_2[3572]) begin
            regVec_3572 <= _zz_regVec_0_1;
          end
          if(_zz_2[3573]) begin
            regVec_3573 <= _zz_regVec_0_1;
          end
          if(_zz_2[3574]) begin
            regVec_3574 <= _zz_regVec_0_1;
          end
          if(_zz_2[3575]) begin
            regVec_3575 <= _zz_regVec_0_1;
          end
          if(_zz_2[3576]) begin
            regVec_3576 <= _zz_regVec_0_1;
          end
          if(_zz_2[3577]) begin
            regVec_3577 <= _zz_regVec_0_1;
          end
          if(_zz_2[3578]) begin
            regVec_3578 <= _zz_regVec_0_1;
          end
          if(_zz_2[3579]) begin
            regVec_3579 <= _zz_regVec_0_1;
          end
          if(_zz_2[3580]) begin
            regVec_3580 <= _zz_regVec_0_1;
          end
          if(_zz_2[3581]) begin
            regVec_3581 <= _zz_regVec_0_1;
          end
          if(_zz_2[3582]) begin
            regVec_3582 <= _zz_regVec_0_1;
          end
          if(_zz_2[3583]) begin
            regVec_3583 <= _zz_regVec_0_1;
          end
          if(_zz_2[3584]) begin
            regVec_3584 <= _zz_regVec_0_1;
          end
          if(_zz_2[3585]) begin
            regVec_3585 <= _zz_regVec_0_1;
          end
          if(_zz_2[3586]) begin
            regVec_3586 <= _zz_regVec_0_1;
          end
          if(_zz_2[3587]) begin
            regVec_3587 <= _zz_regVec_0_1;
          end
          if(_zz_2[3588]) begin
            regVec_3588 <= _zz_regVec_0_1;
          end
          if(_zz_2[3589]) begin
            regVec_3589 <= _zz_regVec_0_1;
          end
          if(_zz_2[3590]) begin
            regVec_3590 <= _zz_regVec_0_1;
          end
          if(_zz_2[3591]) begin
            regVec_3591 <= _zz_regVec_0_1;
          end
          if(_zz_2[3592]) begin
            regVec_3592 <= _zz_regVec_0_1;
          end
          if(_zz_2[3593]) begin
            regVec_3593 <= _zz_regVec_0_1;
          end
          if(_zz_2[3594]) begin
            regVec_3594 <= _zz_regVec_0_1;
          end
          if(_zz_2[3595]) begin
            regVec_3595 <= _zz_regVec_0_1;
          end
          if(_zz_2[3596]) begin
            regVec_3596 <= _zz_regVec_0_1;
          end
          if(_zz_2[3597]) begin
            regVec_3597 <= _zz_regVec_0_1;
          end
          if(_zz_2[3598]) begin
            regVec_3598 <= _zz_regVec_0_1;
          end
          if(_zz_2[3599]) begin
            regVec_3599 <= _zz_regVec_0_1;
          end
          if(_zz_2[3600]) begin
            regVec_3600 <= _zz_regVec_0_1;
          end
          if(_zz_2[3601]) begin
            regVec_3601 <= _zz_regVec_0_1;
          end
          if(_zz_2[3602]) begin
            regVec_3602 <= _zz_regVec_0_1;
          end
          if(_zz_2[3603]) begin
            regVec_3603 <= _zz_regVec_0_1;
          end
          if(_zz_2[3604]) begin
            regVec_3604 <= _zz_regVec_0_1;
          end
          if(_zz_2[3605]) begin
            regVec_3605 <= _zz_regVec_0_1;
          end
          if(_zz_2[3606]) begin
            regVec_3606 <= _zz_regVec_0_1;
          end
          if(_zz_2[3607]) begin
            regVec_3607 <= _zz_regVec_0_1;
          end
          if(_zz_2[3608]) begin
            regVec_3608 <= _zz_regVec_0_1;
          end
          if(_zz_2[3609]) begin
            regVec_3609 <= _zz_regVec_0_1;
          end
          if(_zz_2[3610]) begin
            regVec_3610 <= _zz_regVec_0_1;
          end
          if(_zz_2[3611]) begin
            regVec_3611 <= _zz_regVec_0_1;
          end
          if(_zz_2[3612]) begin
            regVec_3612 <= _zz_regVec_0_1;
          end
          if(_zz_2[3613]) begin
            regVec_3613 <= _zz_regVec_0_1;
          end
          if(_zz_2[3614]) begin
            regVec_3614 <= _zz_regVec_0_1;
          end
          if(_zz_2[3615]) begin
            regVec_3615 <= _zz_regVec_0_1;
          end
          if(_zz_2[3616]) begin
            regVec_3616 <= _zz_regVec_0_1;
          end
          if(_zz_2[3617]) begin
            regVec_3617 <= _zz_regVec_0_1;
          end
          if(_zz_2[3618]) begin
            regVec_3618 <= _zz_regVec_0_1;
          end
          if(_zz_2[3619]) begin
            regVec_3619 <= _zz_regVec_0_1;
          end
          if(_zz_2[3620]) begin
            regVec_3620 <= _zz_regVec_0_1;
          end
          if(_zz_2[3621]) begin
            regVec_3621 <= _zz_regVec_0_1;
          end
          if(_zz_2[3622]) begin
            regVec_3622 <= _zz_regVec_0_1;
          end
          if(_zz_2[3623]) begin
            regVec_3623 <= _zz_regVec_0_1;
          end
          if(_zz_2[3624]) begin
            regVec_3624 <= _zz_regVec_0_1;
          end
          if(_zz_2[3625]) begin
            regVec_3625 <= _zz_regVec_0_1;
          end
          if(_zz_2[3626]) begin
            regVec_3626 <= _zz_regVec_0_1;
          end
          if(_zz_2[3627]) begin
            regVec_3627 <= _zz_regVec_0_1;
          end
          if(_zz_2[3628]) begin
            regVec_3628 <= _zz_regVec_0_1;
          end
          if(_zz_2[3629]) begin
            regVec_3629 <= _zz_regVec_0_1;
          end
          if(_zz_2[3630]) begin
            regVec_3630 <= _zz_regVec_0_1;
          end
          if(_zz_2[3631]) begin
            regVec_3631 <= _zz_regVec_0_1;
          end
          if(_zz_2[3632]) begin
            regVec_3632 <= _zz_regVec_0_1;
          end
          if(_zz_2[3633]) begin
            regVec_3633 <= _zz_regVec_0_1;
          end
          if(_zz_2[3634]) begin
            regVec_3634 <= _zz_regVec_0_1;
          end
          if(_zz_2[3635]) begin
            regVec_3635 <= _zz_regVec_0_1;
          end
          if(_zz_2[3636]) begin
            regVec_3636 <= _zz_regVec_0_1;
          end
          if(_zz_2[3637]) begin
            regVec_3637 <= _zz_regVec_0_1;
          end
          if(_zz_2[3638]) begin
            regVec_3638 <= _zz_regVec_0_1;
          end
          if(_zz_2[3639]) begin
            regVec_3639 <= _zz_regVec_0_1;
          end
          if(_zz_2[3640]) begin
            regVec_3640 <= _zz_regVec_0_1;
          end
          if(_zz_2[3641]) begin
            regVec_3641 <= _zz_regVec_0_1;
          end
          if(_zz_2[3642]) begin
            regVec_3642 <= _zz_regVec_0_1;
          end
          if(_zz_2[3643]) begin
            regVec_3643 <= _zz_regVec_0_1;
          end
          if(_zz_2[3644]) begin
            regVec_3644 <= _zz_regVec_0_1;
          end
          if(_zz_2[3645]) begin
            regVec_3645 <= _zz_regVec_0_1;
          end
          if(_zz_2[3646]) begin
            regVec_3646 <= _zz_regVec_0_1;
          end
          if(_zz_2[3647]) begin
            regVec_3647 <= _zz_regVec_0_1;
          end
          if(_zz_2[3648]) begin
            regVec_3648 <= _zz_regVec_0_1;
          end
          if(_zz_2[3649]) begin
            regVec_3649 <= _zz_regVec_0_1;
          end
          if(_zz_2[3650]) begin
            regVec_3650 <= _zz_regVec_0_1;
          end
          if(_zz_2[3651]) begin
            regVec_3651 <= _zz_regVec_0_1;
          end
          if(_zz_2[3652]) begin
            regVec_3652 <= _zz_regVec_0_1;
          end
          if(_zz_2[3653]) begin
            regVec_3653 <= _zz_regVec_0_1;
          end
          if(_zz_2[3654]) begin
            regVec_3654 <= _zz_regVec_0_1;
          end
          if(_zz_2[3655]) begin
            regVec_3655 <= _zz_regVec_0_1;
          end
          if(_zz_2[3656]) begin
            regVec_3656 <= _zz_regVec_0_1;
          end
          if(_zz_2[3657]) begin
            regVec_3657 <= _zz_regVec_0_1;
          end
          if(_zz_2[3658]) begin
            regVec_3658 <= _zz_regVec_0_1;
          end
          if(_zz_2[3659]) begin
            regVec_3659 <= _zz_regVec_0_1;
          end
          if(_zz_2[3660]) begin
            regVec_3660 <= _zz_regVec_0_1;
          end
          if(_zz_2[3661]) begin
            regVec_3661 <= _zz_regVec_0_1;
          end
          if(_zz_2[3662]) begin
            regVec_3662 <= _zz_regVec_0_1;
          end
          if(_zz_2[3663]) begin
            regVec_3663 <= _zz_regVec_0_1;
          end
          if(_zz_2[3664]) begin
            regVec_3664 <= _zz_regVec_0_1;
          end
          if(_zz_2[3665]) begin
            regVec_3665 <= _zz_regVec_0_1;
          end
          if(_zz_2[3666]) begin
            regVec_3666 <= _zz_regVec_0_1;
          end
          if(_zz_2[3667]) begin
            regVec_3667 <= _zz_regVec_0_1;
          end
          if(_zz_2[3668]) begin
            regVec_3668 <= _zz_regVec_0_1;
          end
          if(_zz_2[3669]) begin
            regVec_3669 <= _zz_regVec_0_1;
          end
          if(_zz_2[3670]) begin
            regVec_3670 <= _zz_regVec_0_1;
          end
          if(_zz_2[3671]) begin
            regVec_3671 <= _zz_regVec_0_1;
          end
          if(_zz_2[3672]) begin
            regVec_3672 <= _zz_regVec_0_1;
          end
          if(_zz_2[3673]) begin
            regVec_3673 <= _zz_regVec_0_1;
          end
          if(_zz_2[3674]) begin
            regVec_3674 <= _zz_regVec_0_1;
          end
          if(_zz_2[3675]) begin
            regVec_3675 <= _zz_regVec_0_1;
          end
          if(_zz_2[3676]) begin
            regVec_3676 <= _zz_regVec_0_1;
          end
          if(_zz_2[3677]) begin
            regVec_3677 <= _zz_regVec_0_1;
          end
          if(_zz_2[3678]) begin
            regVec_3678 <= _zz_regVec_0_1;
          end
          if(_zz_2[3679]) begin
            regVec_3679 <= _zz_regVec_0_1;
          end
          if(_zz_2[3680]) begin
            regVec_3680 <= _zz_regVec_0_1;
          end
          if(_zz_2[3681]) begin
            regVec_3681 <= _zz_regVec_0_1;
          end
          if(_zz_2[3682]) begin
            regVec_3682 <= _zz_regVec_0_1;
          end
          if(_zz_2[3683]) begin
            regVec_3683 <= _zz_regVec_0_1;
          end
          if(_zz_2[3684]) begin
            regVec_3684 <= _zz_regVec_0_1;
          end
          if(_zz_2[3685]) begin
            regVec_3685 <= _zz_regVec_0_1;
          end
          if(_zz_2[3686]) begin
            regVec_3686 <= _zz_regVec_0_1;
          end
          if(_zz_2[3687]) begin
            regVec_3687 <= _zz_regVec_0_1;
          end
          if(_zz_2[3688]) begin
            regVec_3688 <= _zz_regVec_0_1;
          end
          if(_zz_2[3689]) begin
            regVec_3689 <= _zz_regVec_0_1;
          end
          if(_zz_2[3690]) begin
            regVec_3690 <= _zz_regVec_0_1;
          end
          if(_zz_2[3691]) begin
            regVec_3691 <= _zz_regVec_0_1;
          end
          if(_zz_2[3692]) begin
            regVec_3692 <= _zz_regVec_0_1;
          end
          if(_zz_2[3693]) begin
            regVec_3693 <= _zz_regVec_0_1;
          end
          if(_zz_2[3694]) begin
            regVec_3694 <= _zz_regVec_0_1;
          end
          if(_zz_2[3695]) begin
            regVec_3695 <= _zz_regVec_0_1;
          end
          if(_zz_2[3696]) begin
            regVec_3696 <= _zz_regVec_0_1;
          end
          if(_zz_2[3697]) begin
            regVec_3697 <= _zz_regVec_0_1;
          end
          if(_zz_2[3698]) begin
            regVec_3698 <= _zz_regVec_0_1;
          end
          if(_zz_2[3699]) begin
            regVec_3699 <= _zz_regVec_0_1;
          end
          if(_zz_2[3700]) begin
            regVec_3700 <= _zz_regVec_0_1;
          end
          if(_zz_2[3701]) begin
            regVec_3701 <= _zz_regVec_0_1;
          end
          if(_zz_2[3702]) begin
            regVec_3702 <= _zz_regVec_0_1;
          end
          if(_zz_2[3703]) begin
            regVec_3703 <= _zz_regVec_0_1;
          end
          if(_zz_2[3704]) begin
            regVec_3704 <= _zz_regVec_0_1;
          end
          if(_zz_2[3705]) begin
            regVec_3705 <= _zz_regVec_0_1;
          end
          if(_zz_2[3706]) begin
            regVec_3706 <= _zz_regVec_0_1;
          end
          if(_zz_2[3707]) begin
            regVec_3707 <= _zz_regVec_0_1;
          end
          if(_zz_2[3708]) begin
            regVec_3708 <= _zz_regVec_0_1;
          end
          if(_zz_2[3709]) begin
            regVec_3709 <= _zz_regVec_0_1;
          end
          if(_zz_2[3710]) begin
            regVec_3710 <= _zz_regVec_0_1;
          end
          if(_zz_2[3711]) begin
            regVec_3711 <= _zz_regVec_0_1;
          end
          if(_zz_2[3712]) begin
            regVec_3712 <= _zz_regVec_0_1;
          end
          if(_zz_2[3713]) begin
            regVec_3713 <= _zz_regVec_0_1;
          end
          if(_zz_2[3714]) begin
            regVec_3714 <= _zz_regVec_0_1;
          end
          if(_zz_2[3715]) begin
            regVec_3715 <= _zz_regVec_0_1;
          end
          if(_zz_2[3716]) begin
            regVec_3716 <= _zz_regVec_0_1;
          end
          if(_zz_2[3717]) begin
            regVec_3717 <= _zz_regVec_0_1;
          end
          if(_zz_2[3718]) begin
            regVec_3718 <= _zz_regVec_0_1;
          end
          if(_zz_2[3719]) begin
            regVec_3719 <= _zz_regVec_0_1;
          end
          if(_zz_2[3720]) begin
            regVec_3720 <= _zz_regVec_0_1;
          end
          if(_zz_2[3721]) begin
            regVec_3721 <= _zz_regVec_0_1;
          end
          if(_zz_2[3722]) begin
            regVec_3722 <= _zz_regVec_0_1;
          end
          if(_zz_2[3723]) begin
            regVec_3723 <= _zz_regVec_0_1;
          end
          if(_zz_2[3724]) begin
            regVec_3724 <= _zz_regVec_0_1;
          end
          if(_zz_2[3725]) begin
            regVec_3725 <= _zz_regVec_0_1;
          end
          if(_zz_2[3726]) begin
            regVec_3726 <= _zz_regVec_0_1;
          end
          if(_zz_2[3727]) begin
            regVec_3727 <= _zz_regVec_0_1;
          end
          if(_zz_2[3728]) begin
            regVec_3728 <= _zz_regVec_0_1;
          end
          if(_zz_2[3729]) begin
            regVec_3729 <= _zz_regVec_0_1;
          end
          if(_zz_2[3730]) begin
            regVec_3730 <= _zz_regVec_0_1;
          end
          if(_zz_2[3731]) begin
            regVec_3731 <= _zz_regVec_0_1;
          end
          if(_zz_2[3732]) begin
            regVec_3732 <= _zz_regVec_0_1;
          end
          if(_zz_2[3733]) begin
            regVec_3733 <= _zz_regVec_0_1;
          end
          if(_zz_2[3734]) begin
            regVec_3734 <= _zz_regVec_0_1;
          end
          if(_zz_2[3735]) begin
            regVec_3735 <= _zz_regVec_0_1;
          end
          if(_zz_2[3736]) begin
            regVec_3736 <= _zz_regVec_0_1;
          end
          if(_zz_2[3737]) begin
            regVec_3737 <= _zz_regVec_0_1;
          end
          if(_zz_2[3738]) begin
            regVec_3738 <= _zz_regVec_0_1;
          end
          if(_zz_2[3739]) begin
            regVec_3739 <= _zz_regVec_0_1;
          end
          if(_zz_2[3740]) begin
            regVec_3740 <= _zz_regVec_0_1;
          end
          if(_zz_2[3741]) begin
            regVec_3741 <= _zz_regVec_0_1;
          end
          if(_zz_2[3742]) begin
            regVec_3742 <= _zz_regVec_0_1;
          end
          if(_zz_2[3743]) begin
            regVec_3743 <= _zz_regVec_0_1;
          end
          if(_zz_2[3744]) begin
            regVec_3744 <= _zz_regVec_0_1;
          end
          if(_zz_2[3745]) begin
            regVec_3745 <= _zz_regVec_0_1;
          end
          if(_zz_2[3746]) begin
            regVec_3746 <= _zz_regVec_0_1;
          end
          if(_zz_2[3747]) begin
            regVec_3747 <= _zz_regVec_0_1;
          end
          if(_zz_2[3748]) begin
            regVec_3748 <= _zz_regVec_0_1;
          end
          if(_zz_2[3749]) begin
            regVec_3749 <= _zz_regVec_0_1;
          end
          if(_zz_2[3750]) begin
            regVec_3750 <= _zz_regVec_0_1;
          end
          if(_zz_2[3751]) begin
            regVec_3751 <= _zz_regVec_0_1;
          end
          if(_zz_2[3752]) begin
            regVec_3752 <= _zz_regVec_0_1;
          end
          if(_zz_2[3753]) begin
            regVec_3753 <= _zz_regVec_0_1;
          end
          if(_zz_2[3754]) begin
            regVec_3754 <= _zz_regVec_0_1;
          end
          if(_zz_2[3755]) begin
            regVec_3755 <= _zz_regVec_0_1;
          end
          if(_zz_2[3756]) begin
            regVec_3756 <= _zz_regVec_0_1;
          end
          if(_zz_2[3757]) begin
            regVec_3757 <= _zz_regVec_0_1;
          end
          if(_zz_2[3758]) begin
            regVec_3758 <= _zz_regVec_0_1;
          end
          if(_zz_2[3759]) begin
            regVec_3759 <= _zz_regVec_0_1;
          end
          if(_zz_2[3760]) begin
            regVec_3760 <= _zz_regVec_0_1;
          end
          if(_zz_2[3761]) begin
            regVec_3761 <= _zz_regVec_0_1;
          end
          if(_zz_2[3762]) begin
            regVec_3762 <= _zz_regVec_0_1;
          end
          if(_zz_2[3763]) begin
            regVec_3763 <= _zz_regVec_0_1;
          end
          if(_zz_2[3764]) begin
            regVec_3764 <= _zz_regVec_0_1;
          end
          if(_zz_2[3765]) begin
            regVec_3765 <= _zz_regVec_0_1;
          end
          if(_zz_2[3766]) begin
            regVec_3766 <= _zz_regVec_0_1;
          end
          if(_zz_2[3767]) begin
            regVec_3767 <= _zz_regVec_0_1;
          end
          if(_zz_2[3768]) begin
            regVec_3768 <= _zz_regVec_0_1;
          end
          if(_zz_2[3769]) begin
            regVec_3769 <= _zz_regVec_0_1;
          end
          if(_zz_2[3770]) begin
            regVec_3770 <= _zz_regVec_0_1;
          end
          if(_zz_2[3771]) begin
            regVec_3771 <= _zz_regVec_0_1;
          end
          if(_zz_2[3772]) begin
            regVec_3772 <= _zz_regVec_0_1;
          end
          if(_zz_2[3773]) begin
            regVec_3773 <= _zz_regVec_0_1;
          end
          if(_zz_2[3774]) begin
            regVec_3774 <= _zz_regVec_0_1;
          end
          if(_zz_2[3775]) begin
            regVec_3775 <= _zz_regVec_0_1;
          end
          if(_zz_2[3776]) begin
            regVec_3776 <= _zz_regVec_0_1;
          end
          if(_zz_2[3777]) begin
            regVec_3777 <= _zz_regVec_0_1;
          end
          if(_zz_2[3778]) begin
            regVec_3778 <= _zz_regVec_0_1;
          end
          if(_zz_2[3779]) begin
            regVec_3779 <= _zz_regVec_0_1;
          end
          if(_zz_2[3780]) begin
            regVec_3780 <= _zz_regVec_0_1;
          end
          if(_zz_2[3781]) begin
            regVec_3781 <= _zz_regVec_0_1;
          end
          if(_zz_2[3782]) begin
            regVec_3782 <= _zz_regVec_0_1;
          end
          if(_zz_2[3783]) begin
            regVec_3783 <= _zz_regVec_0_1;
          end
          if(_zz_2[3784]) begin
            regVec_3784 <= _zz_regVec_0_1;
          end
          if(_zz_2[3785]) begin
            regVec_3785 <= _zz_regVec_0_1;
          end
          if(_zz_2[3786]) begin
            regVec_3786 <= _zz_regVec_0_1;
          end
          if(_zz_2[3787]) begin
            regVec_3787 <= _zz_regVec_0_1;
          end
          if(_zz_2[3788]) begin
            regVec_3788 <= _zz_regVec_0_1;
          end
          if(_zz_2[3789]) begin
            regVec_3789 <= _zz_regVec_0_1;
          end
          if(_zz_2[3790]) begin
            regVec_3790 <= _zz_regVec_0_1;
          end
          if(_zz_2[3791]) begin
            regVec_3791 <= _zz_regVec_0_1;
          end
          if(_zz_2[3792]) begin
            regVec_3792 <= _zz_regVec_0_1;
          end
          if(_zz_2[3793]) begin
            regVec_3793 <= _zz_regVec_0_1;
          end
          if(_zz_2[3794]) begin
            regVec_3794 <= _zz_regVec_0_1;
          end
          if(_zz_2[3795]) begin
            regVec_3795 <= _zz_regVec_0_1;
          end
          if(_zz_2[3796]) begin
            regVec_3796 <= _zz_regVec_0_1;
          end
          if(_zz_2[3797]) begin
            regVec_3797 <= _zz_regVec_0_1;
          end
          if(_zz_2[3798]) begin
            regVec_3798 <= _zz_regVec_0_1;
          end
          if(_zz_2[3799]) begin
            regVec_3799 <= _zz_regVec_0_1;
          end
          if(_zz_2[3800]) begin
            regVec_3800 <= _zz_regVec_0_1;
          end
          if(_zz_2[3801]) begin
            regVec_3801 <= _zz_regVec_0_1;
          end
          if(_zz_2[3802]) begin
            regVec_3802 <= _zz_regVec_0_1;
          end
          if(_zz_2[3803]) begin
            regVec_3803 <= _zz_regVec_0_1;
          end
          if(_zz_2[3804]) begin
            regVec_3804 <= _zz_regVec_0_1;
          end
          if(_zz_2[3805]) begin
            regVec_3805 <= _zz_regVec_0_1;
          end
          if(_zz_2[3806]) begin
            regVec_3806 <= _zz_regVec_0_1;
          end
          if(_zz_2[3807]) begin
            regVec_3807 <= _zz_regVec_0_1;
          end
          if(_zz_2[3808]) begin
            regVec_3808 <= _zz_regVec_0_1;
          end
          if(_zz_2[3809]) begin
            regVec_3809 <= _zz_regVec_0_1;
          end
          if(_zz_2[3810]) begin
            regVec_3810 <= _zz_regVec_0_1;
          end
          if(_zz_2[3811]) begin
            regVec_3811 <= _zz_regVec_0_1;
          end
          if(_zz_2[3812]) begin
            regVec_3812 <= _zz_regVec_0_1;
          end
          if(_zz_2[3813]) begin
            regVec_3813 <= _zz_regVec_0_1;
          end
          if(_zz_2[3814]) begin
            regVec_3814 <= _zz_regVec_0_1;
          end
          if(_zz_2[3815]) begin
            regVec_3815 <= _zz_regVec_0_1;
          end
          if(_zz_2[3816]) begin
            regVec_3816 <= _zz_regVec_0_1;
          end
          if(_zz_2[3817]) begin
            regVec_3817 <= _zz_regVec_0_1;
          end
          if(_zz_2[3818]) begin
            regVec_3818 <= _zz_regVec_0_1;
          end
          if(_zz_2[3819]) begin
            regVec_3819 <= _zz_regVec_0_1;
          end
          if(_zz_2[3820]) begin
            regVec_3820 <= _zz_regVec_0_1;
          end
          if(_zz_2[3821]) begin
            regVec_3821 <= _zz_regVec_0_1;
          end
          if(_zz_2[3822]) begin
            regVec_3822 <= _zz_regVec_0_1;
          end
          if(_zz_2[3823]) begin
            regVec_3823 <= _zz_regVec_0_1;
          end
          if(_zz_2[3824]) begin
            regVec_3824 <= _zz_regVec_0_1;
          end
          if(_zz_2[3825]) begin
            regVec_3825 <= _zz_regVec_0_1;
          end
          if(_zz_2[3826]) begin
            regVec_3826 <= _zz_regVec_0_1;
          end
          if(_zz_2[3827]) begin
            regVec_3827 <= _zz_regVec_0_1;
          end
          if(_zz_2[3828]) begin
            regVec_3828 <= _zz_regVec_0_1;
          end
          if(_zz_2[3829]) begin
            regVec_3829 <= _zz_regVec_0_1;
          end
          if(_zz_2[3830]) begin
            regVec_3830 <= _zz_regVec_0_1;
          end
          if(_zz_2[3831]) begin
            regVec_3831 <= _zz_regVec_0_1;
          end
          if(_zz_2[3832]) begin
            regVec_3832 <= _zz_regVec_0_1;
          end
          if(_zz_2[3833]) begin
            regVec_3833 <= _zz_regVec_0_1;
          end
          if(_zz_2[3834]) begin
            regVec_3834 <= _zz_regVec_0_1;
          end
          if(_zz_2[3835]) begin
            regVec_3835 <= _zz_regVec_0_1;
          end
          if(_zz_2[3836]) begin
            regVec_3836 <= _zz_regVec_0_1;
          end
          if(_zz_2[3837]) begin
            regVec_3837 <= _zz_regVec_0_1;
          end
          if(_zz_2[3838]) begin
            regVec_3838 <= _zz_regVec_0_1;
          end
          if(_zz_2[3839]) begin
            regVec_3839 <= _zz_regVec_0_1;
          end
          if(_zz_2[3840]) begin
            regVec_3840 <= _zz_regVec_0_1;
          end
          if(_zz_2[3841]) begin
            regVec_3841 <= _zz_regVec_0_1;
          end
          if(_zz_2[3842]) begin
            regVec_3842 <= _zz_regVec_0_1;
          end
          if(_zz_2[3843]) begin
            regVec_3843 <= _zz_regVec_0_1;
          end
          if(_zz_2[3844]) begin
            regVec_3844 <= _zz_regVec_0_1;
          end
          if(_zz_2[3845]) begin
            regVec_3845 <= _zz_regVec_0_1;
          end
          if(_zz_2[3846]) begin
            regVec_3846 <= _zz_regVec_0_1;
          end
          if(_zz_2[3847]) begin
            regVec_3847 <= _zz_regVec_0_1;
          end
          if(_zz_2[3848]) begin
            regVec_3848 <= _zz_regVec_0_1;
          end
          if(_zz_2[3849]) begin
            regVec_3849 <= _zz_regVec_0_1;
          end
          if(_zz_2[3850]) begin
            regVec_3850 <= _zz_regVec_0_1;
          end
          if(_zz_2[3851]) begin
            regVec_3851 <= _zz_regVec_0_1;
          end
          if(_zz_2[3852]) begin
            regVec_3852 <= _zz_regVec_0_1;
          end
          if(_zz_2[3853]) begin
            regVec_3853 <= _zz_regVec_0_1;
          end
          if(_zz_2[3854]) begin
            regVec_3854 <= _zz_regVec_0_1;
          end
          if(_zz_2[3855]) begin
            regVec_3855 <= _zz_regVec_0_1;
          end
          if(_zz_2[3856]) begin
            regVec_3856 <= _zz_regVec_0_1;
          end
          if(_zz_2[3857]) begin
            regVec_3857 <= _zz_regVec_0_1;
          end
          if(_zz_2[3858]) begin
            regVec_3858 <= _zz_regVec_0_1;
          end
          if(_zz_2[3859]) begin
            regVec_3859 <= _zz_regVec_0_1;
          end
          if(_zz_2[3860]) begin
            regVec_3860 <= _zz_regVec_0_1;
          end
          if(_zz_2[3861]) begin
            regVec_3861 <= _zz_regVec_0_1;
          end
          if(_zz_2[3862]) begin
            regVec_3862 <= _zz_regVec_0_1;
          end
          if(_zz_2[3863]) begin
            regVec_3863 <= _zz_regVec_0_1;
          end
          if(_zz_2[3864]) begin
            regVec_3864 <= _zz_regVec_0_1;
          end
          if(_zz_2[3865]) begin
            regVec_3865 <= _zz_regVec_0_1;
          end
          if(_zz_2[3866]) begin
            regVec_3866 <= _zz_regVec_0_1;
          end
          if(_zz_2[3867]) begin
            regVec_3867 <= _zz_regVec_0_1;
          end
          if(_zz_2[3868]) begin
            regVec_3868 <= _zz_regVec_0_1;
          end
          if(_zz_2[3869]) begin
            regVec_3869 <= _zz_regVec_0_1;
          end
          if(_zz_2[3870]) begin
            regVec_3870 <= _zz_regVec_0_1;
          end
          if(_zz_2[3871]) begin
            regVec_3871 <= _zz_regVec_0_1;
          end
          if(_zz_2[3872]) begin
            regVec_3872 <= _zz_regVec_0_1;
          end
          if(_zz_2[3873]) begin
            regVec_3873 <= _zz_regVec_0_1;
          end
          if(_zz_2[3874]) begin
            regVec_3874 <= _zz_regVec_0_1;
          end
          if(_zz_2[3875]) begin
            regVec_3875 <= _zz_regVec_0_1;
          end
          if(_zz_2[3876]) begin
            regVec_3876 <= _zz_regVec_0_1;
          end
          if(_zz_2[3877]) begin
            regVec_3877 <= _zz_regVec_0_1;
          end
          if(_zz_2[3878]) begin
            regVec_3878 <= _zz_regVec_0_1;
          end
          if(_zz_2[3879]) begin
            regVec_3879 <= _zz_regVec_0_1;
          end
          if(_zz_2[3880]) begin
            regVec_3880 <= _zz_regVec_0_1;
          end
          if(_zz_2[3881]) begin
            regVec_3881 <= _zz_regVec_0_1;
          end
          if(_zz_2[3882]) begin
            regVec_3882 <= _zz_regVec_0_1;
          end
          if(_zz_2[3883]) begin
            regVec_3883 <= _zz_regVec_0_1;
          end
          if(_zz_2[3884]) begin
            regVec_3884 <= _zz_regVec_0_1;
          end
          if(_zz_2[3885]) begin
            regVec_3885 <= _zz_regVec_0_1;
          end
          if(_zz_2[3886]) begin
            regVec_3886 <= _zz_regVec_0_1;
          end
          if(_zz_2[3887]) begin
            regVec_3887 <= _zz_regVec_0_1;
          end
          if(_zz_2[3888]) begin
            regVec_3888 <= _zz_regVec_0_1;
          end
          if(_zz_2[3889]) begin
            regVec_3889 <= _zz_regVec_0_1;
          end
          if(_zz_2[3890]) begin
            regVec_3890 <= _zz_regVec_0_1;
          end
          if(_zz_2[3891]) begin
            regVec_3891 <= _zz_regVec_0_1;
          end
          if(_zz_2[3892]) begin
            regVec_3892 <= _zz_regVec_0_1;
          end
          if(_zz_2[3893]) begin
            regVec_3893 <= _zz_regVec_0_1;
          end
          if(_zz_2[3894]) begin
            regVec_3894 <= _zz_regVec_0_1;
          end
          if(_zz_2[3895]) begin
            regVec_3895 <= _zz_regVec_0_1;
          end
          if(_zz_2[3896]) begin
            regVec_3896 <= _zz_regVec_0_1;
          end
          if(_zz_2[3897]) begin
            regVec_3897 <= _zz_regVec_0_1;
          end
          if(_zz_2[3898]) begin
            regVec_3898 <= _zz_regVec_0_1;
          end
          if(_zz_2[3899]) begin
            regVec_3899 <= _zz_regVec_0_1;
          end
          if(_zz_2[3900]) begin
            regVec_3900 <= _zz_regVec_0_1;
          end
          if(_zz_2[3901]) begin
            regVec_3901 <= _zz_regVec_0_1;
          end
          if(_zz_2[3902]) begin
            regVec_3902 <= _zz_regVec_0_1;
          end
          if(_zz_2[3903]) begin
            regVec_3903 <= _zz_regVec_0_1;
          end
          if(_zz_2[3904]) begin
            regVec_3904 <= _zz_regVec_0_1;
          end
          if(_zz_2[3905]) begin
            regVec_3905 <= _zz_regVec_0_1;
          end
          if(_zz_2[3906]) begin
            regVec_3906 <= _zz_regVec_0_1;
          end
          if(_zz_2[3907]) begin
            regVec_3907 <= _zz_regVec_0_1;
          end
          if(_zz_2[3908]) begin
            regVec_3908 <= _zz_regVec_0_1;
          end
          if(_zz_2[3909]) begin
            regVec_3909 <= _zz_regVec_0_1;
          end
          if(_zz_2[3910]) begin
            regVec_3910 <= _zz_regVec_0_1;
          end
          if(_zz_2[3911]) begin
            regVec_3911 <= _zz_regVec_0_1;
          end
          if(_zz_2[3912]) begin
            regVec_3912 <= _zz_regVec_0_1;
          end
          if(_zz_2[3913]) begin
            regVec_3913 <= _zz_regVec_0_1;
          end
          if(_zz_2[3914]) begin
            regVec_3914 <= _zz_regVec_0_1;
          end
          if(_zz_2[3915]) begin
            regVec_3915 <= _zz_regVec_0_1;
          end
          if(_zz_2[3916]) begin
            regVec_3916 <= _zz_regVec_0_1;
          end
          if(_zz_2[3917]) begin
            regVec_3917 <= _zz_regVec_0_1;
          end
          if(_zz_2[3918]) begin
            regVec_3918 <= _zz_regVec_0_1;
          end
          if(_zz_2[3919]) begin
            regVec_3919 <= _zz_regVec_0_1;
          end
          if(_zz_2[3920]) begin
            regVec_3920 <= _zz_regVec_0_1;
          end
          if(_zz_2[3921]) begin
            regVec_3921 <= _zz_regVec_0_1;
          end
          if(_zz_2[3922]) begin
            regVec_3922 <= _zz_regVec_0_1;
          end
          if(_zz_2[3923]) begin
            regVec_3923 <= _zz_regVec_0_1;
          end
          if(_zz_2[3924]) begin
            regVec_3924 <= _zz_regVec_0_1;
          end
          if(_zz_2[3925]) begin
            regVec_3925 <= _zz_regVec_0_1;
          end
          if(_zz_2[3926]) begin
            regVec_3926 <= _zz_regVec_0_1;
          end
          if(_zz_2[3927]) begin
            regVec_3927 <= _zz_regVec_0_1;
          end
          if(_zz_2[3928]) begin
            regVec_3928 <= _zz_regVec_0_1;
          end
          if(_zz_2[3929]) begin
            regVec_3929 <= _zz_regVec_0_1;
          end
          if(_zz_2[3930]) begin
            regVec_3930 <= _zz_regVec_0_1;
          end
          if(_zz_2[3931]) begin
            regVec_3931 <= _zz_regVec_0_1;
          end
          if(_zz_2[3932]) begin
            regVec_3932 <= _zz_regVec_0_1;
          end
          if(_zz_2[3933]) begin
            regVec_3933 <= _zz_regVec_0_1;
          end
          if(_zz_2[3934]) begin
            regVec_3934 <= _zz_regVec_0_1;
          end
          if(_zz_2[3935]) begin
            regVec_3935 <= _zz_regVec_0_1;
          end
          if(_zz_2[3936]) begin
            regVec_3936 <= _zz_regVec_0_1;
          end
          if(_zz_2[3937]) begin
            regVec_3937 <= _zz_regVec_0_1;
          end
          if(_zz_2[3938]) begin
            regVec_3938 <= _zz_regVec_0_1;
          end
          if(_zz_2[3939]) begin
            regVec_3939 <= _zz_regVec_0_1;
          end
          if(_zz_2[3940]) begin
            regVec_3940 <= _zz_regVec_0_1;
          end
          if(_zz_2[3941]) begin
            regVec_3941 <= _zz_regVec_0_1;
          end
          if(_zz_2[3942]) begin
            regVec_3942 <= _zz_regVec_0_1;
          end
          if(_zz_2[3943]) begin
            regVec_3943 <= _zz_regVec_0_1;
          end
          if(_zz_2[3944]) begin
            regVec_3944 <= _zz_regVec_0_1;
          end
          if(_zz_2[3945]) begin
            regVec_3945 <= _zz_regVec_0_1;
          end
          if(_zz_2[3946]) begin
            regVec_3946 <= _zz_regVec_0_1;
          end
          if(_zz_2[3947]) begin
            regVec_3947 <= _zz_regVec_0_1;
          end
          if(_zz_2[3948]) begin
            regVec_3948 <= _zz_regVec_0_1;
          end
          if(_zz_2[3949]) begin
            regVec_3949 <= _zz_regVec_0_1;
          end
          if(_zz_2[3950]) begin
            regVec_3950 <= _zz_regVec_0_1;
          end
          if(_zz_2[3951]) begin
            regVec_3951 <= _zz_regVec_0_1;
          end
          if(_zz_2[3952]) begin
            regVec_3952 <= _zz_regVec_0_1;
          end
          if(_zz_2[3953]) begin
            regVec_3953 <= _zz_regVec_0_1;
          end
          if(_zz_2[3954]) begin
            regVec_3954 <= _zz_regVec_0_1;
          end
          if(_zz_2[3955]) begin
            regVec_3955 <= _zz_regVec_0_1;
          end
          if(_zz_2[3956]) begin
            regVec_3956 <= _zz_regVec_0_1;
          end
          if(_zz_2[3957]) begin
            regVec_3957 <= _zz_regVec_0_1;
          end
          if(_zz_2[3958]) begin
            regVec_3958 <= _zz_regVec_0_1;
          end
          if(_zz_2[3959]) begin
            regVec_3959 <= _zz_regVec_0_1;
          end
          if(_zz_2[3960]) begin
            regVec_3960 <= _zz_regVec_0_1;
          end
          if(_zz_2[3961]) begin
            regVec_3961 <= _zz_regVec_0_1;
          end
          if(_zz_2[3962]) begin
            regVec_3962 <= _zz_regVec_0_1;
          end
          if(_zz_2[3963]) begin
            regVec_3963 <= _zz_regVec_0_1;
          end
          if(_zz_2[3964]) begin
            regVec_3964 <= _zz_regVec_0_1;
          end
          if(_zz_2[3965]) begin
            regVec_3965 <= _zz_regVec_0_1;
          end
          if(_zz_2[3966]) begin
            regVec_3966 <= _zz_regVec_0_1;
          end
          if(_zz_2[3967]) begin
            regVec_3967 <= _zz_regVec_0_1;
          end
          if(_zz_2[3968]) begin
            regVec_3968 <= _zz_regVec_0_1;
          end
          if(_zz_2[3969]) begin
            regVec_3969 <= _zz_regVec_0_1;
          end
          if(_zz_2[3970]) begin
            regVec_3970 <= _zz_regVec_0_1;
          end
          if(_zz_2[3971]) begin
            regVec_3971 <= _zz_regVec_0_1;
          end
          if(_zz_2[3972]) begin
            regVec_3972 <= _zz_regVec_0_1;
          end
          if(_zz_2[3973]) begin
            regVec_3973 <= _zz_regVec_0_1;
          end
          if(_zz_2[3974]) begin
            regVec_3974 <= _zz_regVec_0_1;
          end
          if(_zz_2[3975]) begin
            regVec_3975 <= _zz_regVec_0_1;
          end
          if(_zz_2[3976]) begin
            regVec_3976 <= _zz_regVec_0_1;
          end
          if(_zz_2[3977]) begin
            regVec_3977 <= _zz_regVec_0_1;
          end
          if(_zz_2[3978]) begin
            regVec_3978 <= _zz_regVec_0_1;
          end
          if(_zz_2[3979]) begin
            regVec_3979 <= _zz_regVec_0_1;
          end
          if(_zz_2[3980]) begin
            regVec_3980 <= _zz_regVec_0_1;
          end
          if(_zz_2[3981]) begin
            regVec_3981 <= _zz_regVec_0_1;
          end
          if(_zz_2[3982]) begin
            regVec_3982 <= _zz_regVec_0_1;
          end
          if(_zz_2[3983]) begin
            regVec_3983 <= _zz_regVec_0_1;
          end
          if(_zz_2[3984]) begin
            regVec_3984 <= _zz_regVec_0_1;
          end
          if(_zz_2[3985]) begin
            regVec_3985 <= _zz_regVec_0_1;
          end
          if(_zz_2[3986]) begin
            regVec_3986 <= _zz_regVec_0_1;
          end
          if(_zz_2[3987]) begin
            regVec_3987 <= _zz_regVec_0_1;
          end
          if(_zz_2[3988]) begin
            regVec_3988 <= _zz_regVec_0_1;
          end
          if(_zz_2[3989]) begin
            regVec_3989 <= _zz_regVec_0_1;
          end
          if(_zz_2[3990]) begin
            regVec_3990 <= _zz_regVec_0_1;
          end
          if(_zz_2[3991]) begin
            regVec_3991 <= _zz_regVec_0_1;
          end
          if(_zz_2[3992]) begin
            regVec_3992 <= _zz_regVec_0_1;
          end
          if(_zz_2[3993]) begin
            regVec_3993 <= _zz_regVec_0_1;
          end
          if(_zz_2[3994]) begin
            regVec_3994 <= _zz_regVec_0_1;
          end
          if(_zz_2[3995]) begin
            regVec_3995 <= _zz_regVec_0_1;
          end
          if(_zz_2[3996]) begin
            regVec_3996 <= _zz_regVec_0_1;
          end
          if(_zz_2[3997]) begin
            regVec_3997 <= _zz_regVec_0_1;
          end
          if(_zz_2[3998]) begin
            regVec_3998 <= _zz_regVec_0_1;
          end
          if(_zz_2[3999]) begin
            regVec_3999 <= _zz_regVec_0_1;
          end
          if(_zz_2[4000]) begin
            regVec_4000 <= _zz_regVec_0_1;
          end
          if(_zz_2[4001]) begin
            regVec_4001 <= _zz_regVec_0_1;
          end
          if(_zz_2[4002]) begin
            regVec_4002 <= _zz_regVec_0_1;
          end
          if(_zz_2[4003]) begin
            regVec_4003 <= _zz_regVec_0_1;
          end
          if(_zz_2[4004]) begin
            regVec_4004 <= _zz_regVec_0_1;
          end
          if(_zz_2[4005]) begin
            regVec_4005 <= _zz_regVec_0_1;
          end
          if(_zz_2[4006]) begin
            regVec_4006 <= _zz_regVec_0_1;
          end
          if(_zz_2[4007]) begin
            regVec_4007 <= _zz_regVec_0_1;
          end
          if(_zz_2[4008]) begin
            regVec_4008 <= _zz_regVec_0_1;
          end
          if(_zz_2[4009]) begin
            regVec_4009 <= _zz_regVec_0_1;
          end
          if(_zz_2[4010]) begin
            regVec_4010 <= _zz_regVec_0_1;
          end
          if(_zz_2[4011]) begin
            regVec_4011 <= _zz_regVec_0_1;
          end
          if(_zz_2[4012]) begin
            regVec_4012 <= _zz_regVec_0_1;
          end
          if(_zz_2[4013]) begin
            regVec_4013 <= _zz_regVec_0_1;
          end
          if(_zz_2[4014]) begin
            regVec_4014 <= _zz_regVec_0_1;
          end
          if(_zz_2[4015]) begin
            regVec_4015 <= _zz_regVec_0_1;
          end
          if(_zz_2[4016]) begin
            regVec_4016 <= _zz_regVec_0_1;
          end
          if(_zz_2[4017]) begin
            regVec_4017 <= _zz_regVec_0_1;
          end
          if(_zz_2[4018]) begin
            regVec_4018 <= _zz_regVec_0_1;
          end
          if(_zz_2[4019]) begin
            regVec_4019 <= _zz_regVec_0_1;
          end
          if(_zz_2[4020]) begin
            regVec_4020 <= _zz_regVec_0_1;
          end
          if(_zz_2[4021]) begin
            regVec_4021 <= _zz_regVec_0_1;
          end
          if(_zz_2[4022]) begin
            regVec_4022 <= _zz_regVec_0_1;
          end
          if(_zz_2[4023]) begin
            regVec_4023 <= _zz_regVec_0_1;
          end
          if(_zz_2[4024]) begin
            regVec_4024 <= _zz_regVec_0_1;
          end
          if(_zz_2[4025]) begin
            regVec_4025 <= _zz_regVec_0_1;
          end
          if(_zz_2[4026]) begin
            regVec_4026 <= _zz_regVec_0_1;
          end
          if(_zz_2[4027]) begin
            regVec_4027 <= _zz_regVec_0_1;
          end
          if(_zz_2[4028]) begin
            regVec_4028 <= _zz_regVec_0_1;
          end
          if(_zz_2[4029]) begin
            regVec_4029 <= _zz_regVec_0_1;
          end
          if(_zz_2[4030]) begin
            regVec_4030 <= _zz_regVec_0_1;
          end
          if(_zz_2[4031]) begin
            regVec_4031 <= _zz_regVec_0_1;
          end
          if(_zz_2[4032]) begin
            regVec_4032 <= _zz_regVec_0_1;
          end
          if(_zz_2[4033]) begin
            regVec_4033 <= _zz_regVec_0_1;
          end
          if(_zz_2[4034]) begin
            regVec_4034 <= _zz_regVec_0_1;
          end
          if(_zz_2[4035]) begin
            regVec_4035 <= _zz_regVec_0_1;
          end
          if(_zz_2[4036]) begin
            regVec_4036 <= _zz_regVec_0_1;
          end
          if(_zz_2[4037]) begin
            regVec_4037 <= _zz_regVec_0_1;
          end
          if(_zz_2[4038]) begin
            regVec_4038 <= _zz_regVec_0_1;
          end
          if(_zz_2[4039]) begin
            regVec_4039 <= _zz_regVec_0_1;
          end
          if(_zz_2[4040]) begin
            regVec_4040 <= _zz_regVec_0_1;
          end
          if(_zz_2[4041]) begin
            regVec_4041 <= _zz_regVec_0_1;
          end
          if(_zz_2[4042]) begin
            regVec_4042 <= _zz_regVec_0_1;
          end
          if(_zz_2[4043]) begin
            regVec_4043 <= _zz_regVec_0_1;
          end
          if(_zz_2[4044]) begin
            regVec_4044 <= _zz_regVec_0_1;
          end
          if(_zz_2[4045]) begin
            regVec_4045 <= _zz_regVec_0_1;
          end
          if(_zz_2[4046]) begin
            regVec_4046 <= _zz_regVec_0_1;
          end
          if(_zz_2[4047]) begin
            regVec_4047 <= _zz_regVec_0_1;
          end
          if(_zz_2[4048]) begin
            regVec_4048 <= _zz_regVec_0_1;
          end
          if(_zz_2[4049]) begin
            regVec_4049 <= _zz_regVec_0_1;
          end
          if(_zz_2[4050]) begin
            regVec_4050 <= _zz_regVec_0_1;
          end
          if(_zz_2[4051]) begin
            regVec_4051 <= _zz_regVec_0_1;
          end
          if(_zz_2[4052]) begin
            regVec_4052 <= _zz_regVec_0_1;
          end
          if(_zz_2[4053]) begin
            regVec_4053 <= _zz_regVec_0_1;
          end
          if(_zz_2[4054]) begin
            regVec_4054 <= _zz_regVec_0_1;
          end
          if(_zz_2[4055]) begin
            regVec_4055 <= _zz_regVec_0_1;
          end
          if(_zz_2[4056]) begin
            regVec_4056 <= _zz_regVec_0_1;
          end
          if(_zz_2[4057]) begin
            regVec_4057 <= _zz_regVec_0_1;
          end
          if(_zz_2[4058]) begin
            regVec_4058 <= _zz_regVec_0_1;
          end
          if(_zz_2[4059]) begin
            regVec_4059 <= _zz_regVec_0_1;
          end
          if(_zz_2[4060]) begin
            regVec_4060 <= _zz_regVec_0_1;
          end
          if(_zz_2[4061]) begin
            regVec_4061 <= _zz_regVec_0_1;
          end
          if(_zz_2[4062]) begin
            regVec_4062 <= _zz_regVec_0_1;
          end
          if(_zz_2[4063]) begin
            regVec_4063 <= _zz_regVec_0_1;
          end
          if(_zz_2[4064]) begin
            regVec_4064 <= _zz_regVec_0_1;
          end
          if(_zz_2[4065]) begin
            regVec_4065 <= _zz_regVec_0_1;
          end
          if(_zz_2[4066]) begin
            regVec_4066 <= _zz_regVec_0_1;
          end
          if(_zz_2[4067]) begin
            regVec_4067 <= _zz_regVec_0_1;
          end
          if(_zz_2[4068]) begin
            regVec_4068 <= _zz_regVec_0_1;
          end
          if(_zz_2[4069]) begin
            regVec_4069 <= _zz_regVec_0_1;
          end
          if(_zz_2[4070]) begin
            regVec_4070 <= _zz_regVec_0_1;
          end
          if(_zz_2[4071]) begin
            regVec_4071 <= _zz_regVec_0_1;
          end
          if(_zz_2[4072]) begin
            regVec_4072 <= _zz_regVec_0_1;
          end
          if(_zz_2[4073]) begin
            regVec_4073 <= _zz_regVec_0_1;
          end
          if(_zz_2[4074]) begin
            regVec_4074 <= _zz_regVec_0_1;
          end
          if(_zz_2[4075]) begin
            regVec_4075 <= _zz_regVec_0_1;
          end
          if(_zz_2[4076]) begin
            regVec_4076 <= _zz_regVec_0_1;
          end
          if(_zz_2[4077]) begin
            regVec_4077 <= _zz_regVec_0_1;
          end
          if(_zz_2[4078]) begin
            regVec_4078 <= _zz_regVec_0_1;
          end
          if(_zz_2[4079]) begin
            regVec_4079 <= _zz_regVec_0_1;
          end
          if(_zz_2[4080]) begin
            regVec_4080 <= _zz_regVec_0_1;
          end
          if(_zz_2[4081]) begin
            regVec_4081 <= _zz_regVec_0_1;
          end
          if(_zz_2[4082]) begin
            regVec_4082 <= _zz_regVec_0_1;
          end
          if(_zz_2[4083]) begin
            regVec_4083 <= _zz_regVec_0_1;
          end
          if(_zz_2[4084]) begin
            regVec_4084 <= _zz_regVec_0_1;
          end
          if(_zz_2[4085]) begin
            regVec_4085 <= _zz_regVec_0_1;
          end
          if(_zz_2[4086]) begin
            regVec_4086 <= _zz_regVec_0_1;
          end
          if(_zz_2[4087]) begin
            regVec_4087 <= _zz_regVec_0_1;
          end
          if(_zz_2[4088]) begin
            regVec_4088 <= _zz_regVec_0_1;
          end
          if(_zz_2[4089]) begin
            regVec_4089 <= _zz_regVec_0_1;
          end
          if(_zz_2[4090]) begin
            regVec_4090 <= _zz_regVec_0_1;
          end
          if(_zz_2[4091]) begin
            regVec_4091 <= _zz_regVec_0_1;
          end
          if(_zz_2[4092]) begin
            regVec_4092 <= _zz_regVec_0_1;
          end
          if(_zz_2[4093]) begin
            regVec_4093 <= _zz_regVec_0_1;
          end
          if(_zz_2[4094]) begin
            regVec_4094 <= _zz_regVec_0_1;
          end
          if(_zz_2[4095]) begin
            regVec_4095 <= _zz_regVec_0_1;
          end
        end
        regAwAddr <= Axi4Incr_result;
      end
      if(when_Axi4_transmission_l128) begin
        writeSuccess <= 1'b1;
      end
      if(when_Axi4_transmission_l132) begin
        writeSuccess <= 1'b0;
      end
      if(when_Axi4_transmission_l138) begin
        updataAr <= 1'b0;
      end else begin
        if(when_Axi4_transmission_l140) begin
          updataAr <= 1'b1;
        end
      end
      if(when_Axi4_transmission_l144) begin
        regArAddr <= _zz_regArAddr[11 : 0];
        regArId <= axiSignal_ar_payload_id;
        regArRegion <= axiSignal_ar_payload_region;
        regArLen <= axiSignal_ar_payload_len;
        regArSize <= axiSignal_ar_payload_size;
        regArBrust <= axiSignal_ar_payload_burst;
        regArLock <= axiSignal_ar_payload_lock;
        regArCache <= axiSignal_ar_payload_cache;
        regArQos <= axiSignal_ar_payload_qos;
        regArUser <= axiSignal_ar_payload_user;
        regArProt <= axiSignal_ar_payload_prot;
      end
      if(when_Axi4_transmission_l171) begin
        regArAddr <= Axi4Incr_result_1;
      end
      if(when_Axi4_transmission_l177) begin
        rFireCounter_value <= 13'h0;
      end
      if(when_Axi4_transmission_l182) begin
        regLast <= 1'b1;
      end else begin
        if(when_Axi4_transmission_l184) begin
          regLast <= 1'b0;
        end
      end
      if(when_Axi4_transmission_l189) begin
        AwArConflict <= 1'b1;
      end else begin
        if(when_Axi4_transmission_l191) begin
          AwArConflict <= 1'b0;
        end
      end
    end
  end


endmodule

//StreamFifo replaced by StreamFifo

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [7:0]    io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [7:0]    io_pop_payload,
  input               io_flush,
  output     [5:0]    io_occupancy,
  output     [5:0]    io_availability,
  input               clk,
  input               reset
);
  reg        [7:0]    _zz_logic_ram_port0;
  wire       [4:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [4:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [4:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [4:0]    logic_pushPtr_valueNext;
  reg        [4:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [4:0]    logic_popPtr_valueNext;
  reg        [4:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l955;
  wire       [4:0]    logic_ptrDif;
  reg [7:0] logic_ram [0:31];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {4'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {4'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 5'h1f);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 5'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 5'h1f);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 5'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l955 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 5'h0;
      logic_popPtr_value <= 5'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l955) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
